

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TJQTNYMSYmKvwBqf6dQ1fKQTaCbXWwIZ2i0Qj/xsPBl7jwX0aGzVO1io82n7JrSY/vd49memM5y5
XpgGRs/4hg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LVVyAF5wv2/mnwp8wasr0jrq7FzFOwX+nlCjYuJ9soR1ODNgTWqyqGQdMKcUeOO+xlMAOBCPUL5k
cuvJ7hhJif23EQWvvU26e62cs30hOBBb7aQtA6bgLbucFp8SD+fVMctTZeOb8yLHB6/SBVh+f6Oe
MQvnR3wy5JV2fVLxon4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AM2TI+iZ+NXoK3+XyMb5UQzjUkoo0JbdACL18eHUkvoYfSa1nRewIoCpGG0ShIvR2ubj0OttYGU0
CltqoR7OcEz7gBV33sfaG/Z4IqqugTQ9RnkuRRZ9iR+2EEoK33zGEfZTprRYPPicHxLS2eztEcwL
NPbM0+RJWXaDzKdio8JjstBy9RMkbcI8QqUwWcSKm+xiga8rG9Fhe3mXohfTfksNgnh+5NrDW3Bx
gY49V1+tpB8R89/dXQJNzHD5p/wz+a82idauBEq/AaeHsF+aa/cUncsfAF+NMXM+hZubWs3TABMB
6mnSWOvD5H8qYKodLhoNnrsEBTX00YVMA+nr0w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E1QER6K/8iMRZtejImJPAPIlubOLvRZopcDd3KW58JjEqvfvDS8BBm4BgA5MhsBIf4Dn7HNZ12wv
T42m5fnQW8OVletWvvSD4zPTQQvWkyj0Qph0hfcckswSYUjrElwfAUiAS0eTSI+Wgg/hpFZfB/LT
wJox6umBnylQOiMdT4XS8IoHWErKMhW0S25bTt2hxjZUWO9QUDHA1DeTbYZJsulhsMNpXLxsyCmQ
rYe51/Niqljnu9XTmXln87/wEBu9loxzz0jer0lTV7USPCSgGDKJ11G5lGen1hB46OpDgh8mZ2zM
1hfbeHmjrGZ0yKyUgA4qoZ39Awm5WTJIzED9ag==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Prl2jkWQfvlhA2g2haD2gnOMWKrQNI6iIZv4g/aXBlw93vGOLql1bmdswgcvWE52WQvp7EjENIf2
1YvvpK05o8+n0fq8ZNQf5aoOX95uLwTTv10B3y17I4Ryl088tlQaCO2PtASIhIvuJ3Q8dM4pD3nk
NcmzV4xbagXRy1TuksP52Of+bkAkvhqtRCTZdIIcSUisSsxc4eTMGtNwhBKzTC/T4Q+C37fKKLRe
Eg/hJ8YSR07kr0xSa1lr1/8BMoU7Bq9vTzmtznVaY2YZ9HdXA3RzO+QU4BWOMf977eDYNb2aU5jK
YpHveAFPyOWa2xr7b0YTW4mEjnoNXMae0HLn3g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J2gPaxXXrpwBHNe/SBeuErH5OgTnzT5/vXIB6JfqcPK/kQ++muv+FLBDW/KoueODO2Ww6jXBt5uX
6NBVXxng/boA2NbGiPugsgHJGGCGCa9uWOzr5tYNmpbZAP0rLOgLf9tWbav9Gx/1oO5/TJ0K9ISU
4NEtw81V5ogYG2eB1lM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sFePsMnUWKK+h2p99bZmsUCP2UIq6vID9ipdGEE1PrIJegr7fJPeOggnc7n0W5GO7aF4X+IkQcbZ
k35+ppiurKbtphlbJw2Tm++0qV4GPVoCwpdTbXFU3xnIcHqCT6sZI32QdZCUoMed63tQLlh+CXSp
3t/nuDUBafG+QETpl8oOqZyuXk6iqZslFmm78EpgWxd1l9QaupQpVdIYLA52YRemxS3GJCq0/Hvw
Jty5dQRZYWVg6jsw2m5S8j+7m9yViEhjBFb6CJxXbQQj3iMNY1y9166zCipq03mqFq7VSSHOwyFN
00JiWtlYmkwaQ0kjBxyGiOihYSKrLqCZfeGc4A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 327264)
`protect data_block
vpq0XE/JUwkFZLKlQFurYYiDCiSq+amUeCbXYhSysL6iXM+FLgB17a2kesbne56FQqRdjLojYNVJ
5FWVwSZregwd6w4erWA5oQmRvdu+hLcMWPjynabmPJPrUBh4HqmskEBxk1haZzgDjL7HGFAM3DKE
h5VMBNn7JLZK/9AEs+Ve1LE5Mp3K7sRkxAEOZOAhIJIuicAbQTN5xWq6aSAOrxJfp/n2qky+qSp4
CvK+oMiKsyngh0ehGV4p+Lem24THWWNnFnBLWjiqfoirazbRHylhFOh93cucAv+mzoQEz3Erzoxv
4pfY+Nk27UCj5VKaQegfb02N0bB8dPIunWISwnnlf6fBowDarEuBWPLP5JbcfajcWbumnb7ZWv6s
1gfcpuxCcVwQ5qx0DIAwSunvIB+Y93p3tGyRk4L/3eGI++80Kq09BAipiQ/OThJwmkCHKWvvs3/b
l7C00n7O0yNA1Zo8jf6rJ6ndEC1XzwIZL1G87jZ2Xd5N2hXfqKcWrn6atBPIqWSeYQ4nDqMQtX61
RhubwysLfNhM3o9ENaPkzYJElI2YZfn76gyCqcqaVUOXFm5raIvigRDMbkAqJdK1NRA4JzZttXiH
TV/Fh0U9NLC72z11lphmxhqpm5uPkqbQqlJ15jrL2bNyCdmj/vMogZvK8RJA3eBccBVyUVaoNMVo
KotiCAH8VZju7pT1DvJ6FWmJX8XwLy9TpKMGwLwQ82UL0IKyi7CPWAokRS5LQUEHFyodCV7KnMA8
rA3Sld1lUFuWvRoeNw+dYCO1brVKW7KbOeyi66bL//BVr3grwb/yYzUNudu5QuyuG8gwE86CqU/4
3f+eic5bdk95dR3dZqSLV26/ptrYtNIN79wHO5YM5x/CQFsopiGY7mDJFtzFAHUWY91RQ6BMinDO
LtGN96licLQZzPhgyqZS9ap0zYxEirQWOSFTN60TFFylMocZNy+IAlMU5Iga+jj02EPOhWONe6zC
xapaH7hcKs3YKFjmabsUggsVMs4OH+dC1Od22Rz6X3nSBIJQ0fXxX55HpfVNjcjRgGaSWUuYjOxv
oV/ew/7B1gIoQ2s5xP1TInYukWHgFOs/hJiQoghGx50CqocyOyR8Gr7YsuLXDFG4hKBJ5tbPyYuk
/PEer3cHt0HwUDVGKXEPDAJh17iA1bsE1ZxCBIkoP2WWdtiw1NvFtFlHgR67tFgy3EaZ+VwbSaeO
o8nRHVUhIIhOJblGPSGwOEhOtGIpGf6/F4dF3I50JA7bfERycxvSC61RH+kkBFJ3g8r+TGecvHV0
4rGlAHpsAJk8tUxSFjUEnpohoExt6lO9Fs+w4dmnuXFEnlcrFDyvW3Jlmv29zIi4mnh4zeX9fkNi
6IWRzrXHt7ZQcr8fKwiDvjaVIoSFAYBnAiBQycxZcYaLJjxcBhS0vle421yTQGuWxcNpdTRUVTFh
G6/GFWLzAIOUHNREdlZ4uQ+IBEvL2hT+So/heswspmp+HQZkKIQVHw3kuMj/gCC5z34tZgoCqCUh
VcU/3aoVU39YsR1n8nqZav0WlQjaJrVs6D5gIvwEhC9tA6JLidhg0tRZCzPVvACXwmG+x6LV88VR
pY9evAsfdJBTrsg4LoQDMRijGQZvJOJuQlIvQuUYSkhkWo3WnCloBajSPTaAqZW5jUVi3PiV95Lj
g7bw+l+KwLBXBJT+26oCujVaLE1sFEQyjICX3W+zAjpGa4AjNFcC/QMLHkYBHFjeccGmYEHcGZrC
DYZESl1CsBN6f9jl35gBTb+oYYAG8LzKDMaxd/f2wNmusuvI9aparp3tvfDyqpxu6mQe6HfCtdfS
lyWiBU5cWmAwTfV2BpqjkTub3bbNUKq0W3TIP+lgiJ0WNcQgy3PYHWGSj04AvpXHI0TKgBzqgvtJ
xclKtx1D9zVYVD40oWvQFTjaLvGP+68Ex1nMgrRWg0eqPQlW0ZKYVdGGdF7M0osDQjm+1d64/rsi
rfw+NFefwetrZOTFgr3IM7w3vAdX0+TZ/VDOUsnTdJc2kyW4gBIgQPLyjb/0QFvMOKzZ99JCgIc4
5zWmQq/dicgHpaQmYqs8o+Re1X9OYvd2gRKrM/UGy1EhrMCx6zNjfFa3z/gXb8/fSqNgH+nNcKBS
rukEeNtf6nmdBnLuZojpNAQgIhO8u7dxjJsuVIqd4kuMGLdF5zOjO1faXzgh0ZAx13HKRCE/75OL
+bZXJnNnDYVuweENrAa2uyhJOBfattzXAPxI36TwJk9XA/rhr+oiQ7bEqlrhD+BKGBC4iIxgl9Aq
6uEMlnsQGwP9EzdU6Q801nmlzGjA4bSXTLRrn+jHsZdzKH00rH/58aJV8ZW04dofRL1z5yqDQQtW
LCiDJnQQQ34Jc4UCQaPJD1jbxko2BE5p3OAA2DMaRsxQNNN4juRvg3COh8Hqcq2QAIDx4yyPRU9/
BCi2p6H7NqD265U4piye8OYw9/ZTnCcE2Y2jByvrMwxmqghYWZGm2xtsvSBvZI7MsnolqnP/DQK6
Yr19BjWNwKRnu4heQtc2SNy1TvNhfR5/2iMVkdPHsKyKqpjm9zAP20fV+unUZmoR0elUYRSEwcsa
3BwjuCaHnvUdfu2IsBZxuVch6RLq3aYtUiyrSuhpxUENjMOLMH6cruED75nzA6fXZ/CdezAqwyVI
TfKgdfboEhrEsItKINj+XfPwtw6VmYQKn8Nu0CrYDlIPrsHsDajerH6mTbznXDLmLw9ku61DJ40i
5xrw3UfM5aEJ1V9m1bLhVCPEDhMK82CNk0d5zVy7k9Xyfg8gKzn0IenwPBwS/bI8Cci8gSCyjROe
Jm86Agw2ubV61YkEZT6LUrDQYgml/OoKEZvOdx5dfxE8kaLFy1OEy0QNlsoti139af1qrNTbiR20
+JL9g792Mmg+rvItaeXkMxr97VjYlplkmITPNSxDAeigoTGwTU8Fr8Pkc/v8rif2J0NIJ7nVzeAq
c9dfHie72nS3xaBoZbxjaV3jH5tgVXRt++7dZZRg2DExZf4ehL6XWnTMgxButs4h8siByyV/Tc8g
2xKYeDbwkcMUQRv1tUhmrj9VN08VUZKQ8UyCXI/FTnIkG2kP/nqIxurHV803ef9kPicza5qc09gm
kLspk9dfgxlrb9ku4pr97+bMQSC7rNfTBJP//kFxvKl2DEVECavFjQcCgutXzRm8Mg+pend/bdTh
0dzLhswxGmCUc37QDYHOPZ8QYyx3yMz66tTC1sZnFJlpTKY8Ve5PrsZE9dNRz1Dw7y9BHzi8UTuU
ua/hlQ8YIFjOqtSx1igPFhWTFILmh05F4ZCh+bg1Rir43mwLrngxLFQZPgv+WzdWK+rXr8xVme0G
x0TTMk93gFNfk8CiLcSzu5CVHpQAEO8FxlU0VL4F9S14b3ScVY+8x/0ioLzMZj4SJz3kYI3bA2zX
jSybO7njzaoO9xgbNG+aakKzDrSphpS2MulYLWOkrxL0eOzndngExiP7wColSD2PdL4znNG44EY6
0gQ2M08OT3xH/fRH7wZbvNas/j/ptpQKwRYeYprzpniu8huDz7RCoKm0w3ri7m4rCAihFJiMSqpf
NBOUCL8WcFXCrzrYkBIEGur+erWIU60KWFaGaFkZZf0I+ilGtvvAU37zhgmoOxQ6fCpFCke7B6hJ
mHkLYh2u1ez4hnKEGgC+3Y0PuwIUwm4CtSyYZhogCn+3GcXOlFqLVrkOfdsiRziiXcT44gqJr+Uc
IcD8S/LCR34aDBPCJpkQO9FYV053WAu7irAPHg9ueuFJFOt7vV4nXzy1efIXlbgWkUIxCooTzpSn
Eqo9erZeCSh9srCg/tQvrYWpfPo0V+x63EuuSvB07s1g0T7eWZUeyiusLg8tOdpmjJspZvIByAaD
1Zb+ismV4SzvRHE+IhFf5uE9eHS6wxlSXn4wFoQGbLMVNQCcLhIuXBj0ZFmIXr3l4C+sQSvM603t
FTHNlAz9Cy9lVUdDQ7nfxwL6svhVFB8Y5fGZtfqWB6jAOYL2w0tNja0bGddYZXLgSEiOhZo3Foha
GnMY+f8WguvlTplp1yGFY3DD321H3MrhWg2vuAixvHnJIDnLZZeGENTfKIoOL68h4nyg2REUtHZF
ibU4qv0alw6HZeYDIfLadRsaKNyuaIUlnroI2t/6r7gi+9MNFGK+TAFPOZt58WKBtwYfCWD5bFvD
p/85opbSAOIYFolTPQMs3s65K4BWB91QajaGCVD9bwNzVqo/e/uM7H4ZZLMDYe+L+Q527SzhJBSP
u3rf6FPSFecpo1Q93K9uabuXGCDdRfSGezprBblzLKvNmfW+vArtzBgHLDxQW35pHpeXHehdH5t0
HfZW8SOBERD2mjbo7iUb3l62PKhAueJmJxjBwhVPy6nu7vvYZD6sQOAnbb1IKa2WHwnIWyya0/zS
3h4az1PdplT3+d1/fjycoRn1NLTfLtAfkuSd+yPECLN8l2WuHuT4JhpVbhJ387tQLIU/1AIV4tHH
D1eWqXjCBrqNqWgfzfSzMiHKQwzPqQCHJ6UxDj3ON8qLsXtsU3mfBqQPoX09iHFyJP7LJw7ZgCAH
TD+n+Xcv6aUcbxHsbzEXf7odf17iPivKn3+UvLQ5En68tKunrpTVdvg19Djajj/O5xTsLM4LhXc+
vu+POugndHJKvVn1R0nNsSZxSU6PjEg+hUahRZlq4e4L1TC1jxevZT84eS+IfwiiqGhc40i/Ssm2
ccR/z3lVSE/K3sR5lr8ZdRNOuTWC0zdgbXhnq2oiiRWv1FJTzqon9z8AYSRjE6E0QtEhvX/Z/pR2
Mg8dpRRHnO0Vl4W0qyI+jpZHe0/ItW8SNScNXi8lrvpLJMAIHMiQX0/LFb5Qbjcg293SS3l4KN14
aaigPGLl8s2L+LVeBpLBwVDOLCDr2hxbCx7uHjy4NXhga1MC9ieEmYA/Nw+ephRjExD/9ecNVple
v0ikTlWLxOgv/dw7gPa6PBCUJNBpwl6m1tqcEBK60jdsTded2l8b512Bkt/9DOgmz5GKEt91xFLu
1sWg9E1Wojy1EYlfRxavISZgVrEN/ZvC2jQj5BN16w5E03IEYXfCC4Lmv9cddOEZW8B99nIzjRRz
QGixg2kTNcDquUIwmp8mNUBrEGiyn8PBQYjWPUaq0KGXBwVq0R+7Czj8FlrMOXtxu3mtpK2LuO9h
PdtDrOb9xNBH4OWkda+qW6dOXcOyVLpiEwlUWENWAyVNtEuvzbVw2Rp50AB36pvaECrZocyI9u5V
fYGFrV9pYqImmxDFG4SYlPy8Bgl2LZ2XdNn1NjWVEiAgvM2go7t4IMJ+WYPvfrALCvvSX1nEf2a/
lytJs43dd54is8s4mYNZdE4fCs5RsYcL/J9iH9w7M80L5qCU6sL7rwXK31giAnOY6qUJBSCC02Es
N4jTxHEq8vsVYRugW9oyyi0iwRUFu3Cj8R0ioD2O+nqUr2g+PWdH2bHpSfQ/SVRYC1Y4mOHAjSdK
cPEk5B6nDT+h292xETlhNfbqAnPFH5YgmsCRRT/NpxrkkDAvdglS6SCUy6JHqDtPgOE8/RSYya/u
6advkzk4BXhU/E/Fpe5gjTPF7OMLDkRTxIaKCGmUc2IlH/lsnPR5wPin+A063MtPYGJp7O7P0Ls7
UnFC+Zl+yKMuhVG8OhMoyu9Y7xRTTDdk/weHqd3MjAdE/yk/5WS8pADhtmd65GLaxjYWcAZOvZLm
7z85ox0HbpDmIW25sHS/BPy6MSYkAaXLyfd/HXDUJVOwJ6gaiEKN4m5gyz1HS3Qq1ZT52Xh8z12+
K3UXgRf4EbDcuTkYXN6VraegDN/ZcF02MlkJBPug41I5UEizyUNCnhA+5fSJ6WphN3q2fYYSHs4V
y+zuDMy5kbp5HMw5o/CJcbdSTTZpc4cdasWzVfqx7QsDoOSOyZidtEJzC3yurv1t+KbbEcJv8d65
oWWUwmimN+aueP7rM2uw11A6WI3Z5+jnDkb9LCG7zCFAOkrdmx1WUHmdBYGvhopwPtPTO0AKUTWH
jhlz1WsQN/4nCKam5awzuYzgZhKcq0bPiefAFDUslw8wi7pVmbMpFUTdwkaoSX4qR53FdGpkwg+S
SrSdaulB6tA4fgjLnKkAbgA3/MVOmFKHOodNOaCiJShYSE9p8vlfDBa+nseSRRsFHYwZulKvBosW
QctU5H1rzRLmS9uYbSBfCyOrZRt2Hch6/ZZ+elpPmEtCHeWdUTZxlhh2bY3hVgBsm4rhp/ldZStQ
0PJlSeSyJQR78M5OA4xmL+WS5PVPP5Yzgxv4N8tMnKxy9SbeZiuUKsPsf8LvCjS4SdzN8qD5+JXv
gCV1mn2ku8gJWdKr/f5xOwORuEKVulxfrv1O6w0ulUlpjl8fzJ/DprKv+bnDjczIN9hoNifm1tnS
NFacyHNr4ncdn93D00tXeG7/7np/El+UGmRKKUnSMZSrq3RdWejoyZ4fiM/AjCIkBD5bWNM5fyDn
8AAzhtU2o1hCWh65wpHlC1d2awcyoh1Y6fKKOZ2nGop5T/xBjyeDvYGz0fIlrszQ5+ckpbp4i+ng
tk8Tu5udtA7ez9a8IP/qa2n8TX7CrweHcPwxAT8UsEdHn8W6UmMDLO0ybR7SkXReOQTN/yMBgHQr
rqwNTpVQer394otg2jahu2CjO/WKjoC6Bbr/3MxfY4doGwmKmCGLNz1bwPBQnqFjAuxhDd3hdl+9
S1TzoYHK2TUWaBbwgnONMfnGFJWW55RkGJvLGHsM0HbHrrbaJSAGthv4fc2zDCKTVb47l6hvkvXT
OObwQUnQet0pRXuaWG37zq+4QxVkBxbtxOiIFuzeZjoyqBPjy0bnmL0u+ZXuz/AkhpjiCCBgGQiT
WR9uwNZYpJdcNlmTLCnN58KjqbO2AuFmCpegMEWpKAWT6/x7Bj9Rl5EkqUG2Y87n8WUhJ1lgIcXr
FNUnMBpnqjAZt7C1u5z7il3aFlfvmexaTt3DunANWV82+KeB+ggGhzIeGiTyLON6FVbuzuHrn+TM
mL7ZDbJEE6cZBt02AT3zuX17Xn1f58yRvmZ2lvfBBPmCgmqG6zB2aIR1OGBnpsfcPejrUQfE96hs
iJc8XOJGQ9hzh7ErNcHp0FAGZgknWUagyPIWZLzYjWKyFeSKwJec+yzRFi8mSIjAUv0LJizjQ0h0
ZZhZw2b6WrVTi2IR4IFkmO1MoCs2z3j9lXmjwrOpFA0VDmmHwn2s4qG1GHvNWcDI3yD3wsyLoiLI
1CRgFQOAKbbvEi1yUTa624flTfKM2QtGySXBNiKlp9E9oAL8ggic8ZiLmTU/r/4C6t4djRYXvjUr
X0ims18O3nTijgOienaa7RhG+1izwQAYFXWu9zAuTNGptIlnniJ5JnaWq8OgLxsEukLXjPHQjuuI
KTyBrg+TCtIY4jizkY4QbZ96LnA1tFthqFVj4HhAyYfuuvVNewV3hSdc+rbINJ6Dgg/UWDaXRAkG
YJPvWBlJv5KAdz9t+/FLBFVLC4SW+R7M74cVvelRHELHtUysvf/FLJBIOv4Wo7bsrG5nHptV+jOa
fOwXkDqWPzjonuQWuvChcI4q32Qhzyx5GFQmrwh59o2nLnIMmdEYDnlJGtnNe/zcLEVrMnwF4DQR
YYun90SamEf0s7ILIAxQgHgd+K5Zr8ZMw+oMhHzkGc9UENCTAZgRPaPoeaUjhjqsJJZyaXgJziih
IQRwunhAc1HBOmdhB3ocWEzzxazLz6+q3dgffHjck5GtbbQQ9ZrSA5RLTsaQjly8YnR3y6hpTPZ8
/ifizJEb49ycTgfQ2ZwoX72AJ6cugQYICha1AMLlO5xAtwupROKwldVjIyIyLyGgNPyHdxBXUs5y
72DbKZggbtc/oGiWr6Yrs7w6qE5aRfqZDAXujAoCnxHx6myFQC3b3n0SsYNEHH3BzZHTQKAdlluR
F/amGthEoDjMVNmkfJsem5KOfXBtvUrs1Aau5lNg8K/yW7DjH+Kt4cFzj61Lufw22Wesei7p46wr
vRxeGto1jN3/ZjqXZOTN8mNbU1EVpyhmDOEtmBIm41eXhEqrahTjiOb/NG1et+450ay1KgdE5NHq
LnRJiKTx9OJ06vYLy/QcY2j/iDuyvYac4EW6w9pg7MaGi0gXrnv+iKpDEAzYhcksHzmlHi0Y5Oef
c7EuNb87vTCH84fErp+b08e5TtdK1bCDr+FUi+Ir85xXOdr4XXcWYnFbUTD3HKJAlKKCw3MYzyYh
ivLmiPYgWiX95mfvU5p1AHPfFjbG/CtUNTyxXRGZH2Dy9gAVSVjY1VO1BHh8dAapPYrsW0WKKNIx
II8e/3VbyK2dESLbuc+hi5XikmLLSKD5uN/aRysRrMZ8bIDOkN2a/19EwJdVbNhAd7lrl1p97Hx3
331kcy/cFOvEn2QJ7UTysOE1qvbEnmzWEy/h8a0h8qMCW4dN1IWd4Ux1dqbpRm+g/fNO9tJ0Kh+w
yzDFl1/ALX/T0StJ7tMwTfPQlhmNya+P94Aq9wbPdMi69VaykVpMt21WRjzegDbHgxb7ny+Hfcje
rjdzsso5qs7g5t4UFRrSp9tltoZ5aWUJyvT94NrMdFk7NtFaHMzIs9kmFwG+njoWVqD5Pd5mAuPT
jP3uvqT1ni/wdcrITHh3bufFfcNJgagq6lXR5TnVd4jVGFjR3gzYcXkXB9LJ1zz2VRiuyuQCliRm
yQnah9+/dEsAN7JJB/ZGiYKG72qdWCM5S+CegkrQM9movr6DfPGDmPPKd3ONQ8QUgyxOdRHAK/K3
HGwZ+qqSW1X8j/ziyi23WuQpqIFPVJFBH3lKj1Skd2Jket5/gMoGSewBk16fksYZIQy7DGxah/9w
KQzUnhh/CGnJeys4k+c0cmxfa+pc0//E/Md5JfTOcIU3l29rVbCqjyUNJ57pSniI++MOLfFZNUEe
LS8mzNXlaHslXU+ZQ/xZzxLSAgPW1l/ydUm99bBiCqbdcq6WK7su6wfbqyKpHzG3OzqoC4ux91tl
XejTGeXqkn58wlHaoaA0BG6eWrW6PGVj55EioVX5wKWGiGD7him+hQPiUAYbbgtPQ2fuwUGLz8Yh
nhcSdUjyg5Kc6EA7y+UQBaZpAmiawX3BXjPKtlRKHXIvOTswYjXo52qqz+1y9ZCvcwwOKxD2Zq6b
LQlws5dMOQne7AbO6ME3akhuZTqZZZMTn6xp+BWWaDcUJ2J10JCxtQ7pERhgPlJqQxsem6CvicPG
GhtuzVsapzwhJL42sHw/OlvWIlMhy6P2xF99hpp0xHlGvlUOUS4dDTPsB8NAcrsiL5F00dyMsvAA
ghcuS/BzmnlZE5HGusiwHokibSxfaP7jDqQGVkhXa97rpleJaCfd6WJJonCjOSuy+QSM3LT1qq6b
2Nasd1zZOMGPwh54b8a7S/KKO4TDqfCYcisOWTDFkETZh7aYgBbllz6E21IgusyAW0HmA30R3/up
4vej3b58hsW2QQoSuTvDxAkpCH0IBS4CISUk5Z8OFuaYS8FzHC+BQjY8colqmjMZb1yK28OGwQyW
cZFDuhmKmmc3+GWNyAOhOHON/bsRwjYoSqqEviNYXlNMVlxapZ1XH0OJIKEN3o5uNnM49K5opBpz
F701q6SrKVhfMU0CAK+/QySr4kbNBh377wXWvnI61zs7ql2oR6fRh0ypCgAN0uEKM+EXJ1Reu3/2
IhNXMW+EAQ2gTwClNjhFAYMi0olx/mSg58eKI+luolYjr0erTDa8659+Mi3pi0fU1uqz2i8Opjur
ALPnFaeiKu/XvWccA2efYG9FayNBpDNSZM8/qvbVnJXZbjHiyQpIpfUTlVcqxPxtVVI6/GN+vy5A
9jVUujkS/quK4OAl0FjsMnfBRFmudIxoO7puuxrm/abYj6LWi/m6zISJXWX/nAZ17u51cxC3neXu
ibDcp25iyxuU9hFVO593HKmBP2+XrQWmC3pZZoixRQhYqOl1efdhaxtYNn/dchltrmC1BiZElvl0
ZrFS6wNjjWEKk8hU5joX6vA3Dyo5iQ/KMIAazXr+RAuu1BV5F2fpksSpF3y16PNhZ/mDcJxWwjin
ddv410jy9ENbJOsBHjw7icK8jalLfBrA1jJVtUCAHwJgWKk2BblmwxHBEiPT+EoDs0QR286STgV4
7wT7YMUfhB9Rq6VvfBXmDrMOHX5Afq8Ykz606sGTYrCwzUBQCBP8iobgRAy57pK88EN+QKuntFLo
QP/IahJGndZsztVXAoApOjHpltFam2nE5RjFfam6VP53+23VqIB7Q3il+3T9GahVolpEJbNR1zZG
jCsvxUYBcm/DWp59DYR4i6QI5ZCUD9dU3Vam0P9LmA4K+UU8XNuhkP+dC0aD8RozjLQz3542O6hu
NfEIoJoUpL9cFK/g1tvY+kmXXgaobBFjVCKrCaD1+BuDWbVy3iynbmy7qWAO6MUeAeN5HBAneA7j
gSW+Df/OqZf0dPLLkHOXLQNI61WoMfykBaweC4xwEkhSwq39FkECj1kfVkrfXjSaU9QoLZJIb4K4
7h+XxCEHswfXL9ucnGoVOpe/yNYAE6yBh26uV4M+EllIfKPIazTYh8Ib1fa7UZhdRLA6wN9xoo/v
Er5J86nzD8hQ1KwvQ+cmI5RM1eN43/K+Dd2kmcy4P728cwcmHkt2HuXDArfWPy+8FYkJcb/uAqM5
pI+ChMG5hNiGnzPvfKD21EXafeT5Dwx8r1Chl/0+hmqZf7VCBoHVfuW2j0T5vslb0BAuILp6Q8Ck
EroBiYMTyLrY4Swtjw3qKNOKneWDwKi27Uj3dnI3tQjL3i7/hKktAwO51cRQCPtZiY73ZNsTHcba
QKhzck2ajbFsYp1etLyaR/WDkrEWy5gvbLsJPQR5cGedC44JtrpVQhtSdvuGaJNxvj2YOQimz9RM
/VinxglkraOiRmFKe4NhUhwVkgtFl9exWW0jXmGmK5jV1n/CN7IyAYUxDtkXPVoD4GqgrXdKS1L4
7Q7aPoLN4NCQXI0tDS0HFWEhda9fz3GoJ+iVyzD6EmN9Xl+QbCdwNGNiQy9mpETdeEOLbzgJRPAB
Jsc6TEoqCPZoXGJ39VOh4RJaKc+Jt9LlBBlx9Vq9fYvOluToQ0+bCJn2m10r7dTSofYHs+QR/MMk
ebULo90hOlFHzvhj1PVUwWxOYZB2jlpV1HPrMi76NjN+5CN41hGbMXGMwLiKJvGTtDBYvuYr2nIi
0LVcLKTbppnfYD/Nd2FHlZlikhfRAVvz+l9jS+WHiyEQhJWxUQp/vHH6ZfsZKEZqWVhikeFGErLl
tTz7iOh1AnmJNwAQUWMe9tjt1AnOBsVQjFauSyfIsBNDMC0VWYRBl2dZUBudK8yIypi5gcafAgrx
497q82N1H0B4+3o4uoDabRwVY/2xJ4h9zh2vxVBdQs0jrA2lToLtaYNywOZPhC4zo2JC1JxeJaJH
jWrbUEwwnWAMG40Yk9FoS2w3MdUYM3x9Ms6l+orMufC6m4swtCq2SPZABm2XQdst7gR+PQDcYxeY
Lc7fS5513PnVw6/n9D1aFrfkNPCtMDEq1fKWxM+Zk9A9hm5wynLZGwBSwfSWLwGH3OtU5dwVbxKC
ud8m1xSaDyU8COvGU7fPLz/bmhTatCCey45Nq4l+WTQu88g6gWRmt14HjmjbDDJUH+QXydbEBLYS
8Qy4fs/RqvZzC0QVA6bY2WKENaPpc7FWe+QhAgw/GjCjSQCI+cSU+OLDvAhrV5qmeCRrcTOIToua
n72qvWvFMXoEqPnXRIag37jvOFTerj08sfJ6v1ry6eYioYNEEkEZ+FU2IVwk5z/AURT3NmJYkIMP
BzD5VwNnpwjGkV2BDLxOwNnHeMVOMQ+8DQeR5sW42gTiiFlEaactrSJmQGpN4v0gKLt4jlYogmtJ
Rg6yrHZxf0zcXitU3t+FTTTGQNDMuaw4BKJYB9yYRdc0ARejfTGbe7JKoWpZ1TutLZLmC7j0XhLl
hKB+AW0i7s0SBBHdjiMpja1Nm1HR1XqVFHx6mnTiJ1qiM+DRCc33BCBWqVJW9P0MFndk0+gRYSRS
L0UwB6Alzg/VFNlfZ781ICf5KklYOJzMGWs2cAPLUiZQ/gfUBR6Ym7tFVvPxyDfhGl2rMLPcIWAS
tDN7wNykf70gz6eqwQA9uusN1aYywrgZZuLSns4uEU9pSjLuTfgWiqCzLMdMhk9a+pI5m86sREeH
bH5kDmh0iMRGiyXTQdo4mustemanL0LcsPhH83Q6qa6PAweqlOYnC/XdJUd1nIojXqqt+cx1VNpD
6tDjGPtM6OgTWSSTXrUF79Xqsz6KlV70rHmn5R6sbCFNstAM0P9qkwegRjU5DmCRSUe5/+asl0Tb
GUoVmSbOrIyEDC0k7wsynQuOxx+iqCIk74HTvvm3otuLfyNmqjUlwiT8r1iTuNwRz3dIm9Ae5Gqf
4xtNy4dfO/pmUj8/9YgVMGqGNpZOHZZuR0a076yuMnE2LPgkAqLTsJUi8/ZXSHUhFyZb1gzqUT48
xB5dtU+NK6hvnuOh4FBF/upyZ12e55cKzLeozXageeutA4JSkbQS+fhs/p77sUdMFADQE6gxsFpn
2AZNKdKw3bz06t1MygOYax2M743CaMKtYsz6LLi4ycr4MYGPnj1GmKNU6hKMeZG917Nt9KrfMJZo
jz+0f3KMfz7yT0cIKx4s6+aLCMb8nzLvhBax44bfhMTCK6E9DZKProYsF++Bp/ZRQ2VkFrktdgOx
yNCQl8zARBxJvbENM8A8rG7pZnS4RCyGhSK9QfqEhTOCIW6byxywhLAgXQYYVgOqkp0ZDdK/dfFm
rjWA1TyzrxeWBD9WW6UNfyJhJ0KNafOrTc/OI8o72tzWC4tygFaW42ahhCa1AAo38BT3fV581en3
UoBgGRxSYrtfh3QO+0L+x+VyESVS29+zgDm3MvAq82ronP+xatYendqH1ZI78rqSR2nBg7VLNNCl
o4dW0TlpMt1P4t2HKlyQRSpoC80J29re2v4HheEwN1h0mFQZWVRd5IohYd7beuHinYCPCqm1HRuQ
Xn7Jt7OE7XKGk6VadfvfCY/u1R9v3/7NSEUBUdwML33HPHSBSIpq0tzjbPwyKLVTDoa3gF+wQ+z/
KNOiUOxUVX3NB4mNGpzLoOtGrGeaTiCpmthYbgKM1XeS14dNif2xJO1h47HK19nLx1UTxZ4vNewq
+sjDZmyPBKDkg5Aumd7vOgcUWQQImGoZ80QqIO/JUXCuat9NKq2BMkAD1kA8JWP7piRr4kFnyiD9
CKMG2gPTKRRckcKtcccsp5OctzWv62G3doMqlhRU2PgKPB52I+TGlfGrVJTHt8vapfuDCTvKQur7
WV5oHw8zjtiWlEVxm/uD8b0sxnCZHRXWGEb7n/wqZl/mZGBFNzaS1uas/Q5LqE2ntxtXCm4/sKnu
ySHaTZ4PDILsw8hxKrmjn/pg+cZTDUqwZgmJfquvw2AGofbTyDn2of5k2jFuLpx99IRBT0o+1GEu
lIOQraQwLInWlWG0opBRA8uDj1ut0624oENiIolfskE1ysi0Td9o2t6TgQQ9iLQVfFoxSXyqyr0J
3VUBHMazIt/H8C5vvqeJnRwsJFAIWPz+CAiwKWx2/ujdn0t0+7gB/oQDBFcH+pXzNqdrp7VrZBXr
W04LzaRULYvhvbdaAgUlCfuoytNKuOYMFCcD4Ni9mmHK+uF5YEfSTF7LY6DR7xdXy5xdJezy27vu
DhhIdApGCbIiRw5yxeg0q446YY+6SiN1afZQ2bsfJiTQPj3y8R3NzzsxXx5WfUQ+pc69OUAy/fX1
bRl/kbbep1uPxwg9s+cDCWK1wnOx38riOOpNHiiHSNu2CMCBQrW7ixYewV9v4bAWKOcCoTh2w280
Px2s6+457jAGjWysl8Jk8nN0uaj8vCrGTB8A6IkxW8LAWsTLO6/2lKqfNmdmNiwajQO2iSsaMh8/
Wcullgan+ebefeLe9uUpavyytOO4c7wwHWAGu+k/ZlIPwXLTxrOP8i2rjX7D6R+rrMuiA7an5BPz
XjmcUzjhNRZ8Epg5IaLEStbqFGWCfYO1NwrIZKWMocg6Z1uiDfIBcccqdKWvHI27az5lzhgM/w/g
/sTqK3FCLgLhi6RWspbUahNwZNq02t5SjFMkSm/QjnTqbiA2lVyrjQ7yalv/eNPhM0zCmLPaNTeH
CmETLPv7zd5CToQSmauWr6eDIg+6KeTrhCdpJd5dvOgtD039AoFdLfcsgMfrWXTbZCFzwZgoqpBY
XPOhdC32Te2OuBANUPQb6C/yXuytbct+MACKTIQwU9BM2t0pLyQmgiU4lyXK4BkCAM1LaTXBM7p5
V7EXWdMjKziG94EXuf9W547DkalmletwaSijDTbWdXCCcuvEwxEwXke3UzcMms8F4qK3o3fOgSFW
LgcPcPwXxD7mH5Zyrqh22khXC8BeMi5du5P3Z0BdCPYF39l8/kq8d+cAp/VYqMw5Mkry6WYFt0ym
HLExFLHhTZOsmoxP/1VSGIKPsDSdcl94LN5W5TIfxtLZ9tev5R1+Lk0mCiQMQSy9E5q66PUetmEg
Wjxk/MGwwFb/cSnt5MJG+18M4j/GHySlZ7yM3Cz25hGU4UllW02t1ywLtqYMB18tDt6SvmOPkySc
F2AM9xweT9VJGHyRVHg9moLK1CFXCKZrABUv7GW411s/UdBhP3coD+NNOlpIO0XAVLRf3hvb5hD6
UGQ+1x0L+OkaX9SuTIhRviNamAcq6IG4G5iGaBSOig7oRvMUD87glnUUUw26j+8Nk7udZW6s9wR4
WPvWxhSqmCn5aTZi4AmAUgAAW94lxIKwQLX+tzdDKwz+PFqLRZyNdpnLinqAvHut/0VSaW48ZVyX
ydWRrisEL98o0qgAvRCnVxz+apU23ZsJRmoZQ5q0c1iMLAhzFaQSYxMqi0zUnvHPA6juT2jBjKRv
ZsqvEjAw2SU+HoTZSP/aQhhwRqfmN9/bl37uydUIkNkBrNc6Ftz8Jo0Dy8ACd8p31KmxCWZsnHwb
mhAf9tf/W0az/ktYEsDCyIfpMVHhWVUCu2A86DY37z0d3caSX4knvtUqoR7cIyEq+fDSUk7wiRm7
tPxh9nEGYg0dfLAkCe6cHY6jmwiySM9P6v7nIoF1nuzShQt9RSMu8tj7xNq1VMNtQjcp4s4cH9FP
OJKQqPCVANuSfr6tYZXthaHbiXBn6y+MbHm/ZS1voWq2mgjtdCEr8wuTDXjR1BQTMLJj7dKn7p2v
jxSbOcNqqoyGSsl/D229WK2yfgVu6Zul171v2N04J6LI4k4OgMDR5HY2KbnkXC/ixT2saBL/SHLv
iGAihoXFIE0yf4HfyP6xFxXqdD+DLJFs8HW72o/RKZut+ovHwH9zdWPnfj3nrZYf4NlOjKzmZtVw
2Rw4Lyf9pcdWGzkMIZp2DGRPJXeRgCvKAEiJ5D0tydtMSz69CAzz8en95SCVrH10yvxlkXl4sStO
lgeGTJXLKxJihLePkEUcCr9GnnsG1BZ38XHstgasST1QT9sADzO/LeBHvKm0gWF5tXq4TRgOqlSK
VooNCGr+QXyrXOpaW9b7/jp2MH4mXfNTFbPCy0ZiPp/rUQZEca0T05AtjvFKjniK18y5Wdjc6v35
oev5pbEx6AAkHl7PLHlWaSazIhHXlwkkGdjgk0LOimACSXyOixpEatCi9ZZLR20lOpyEY32/rLMC
mU9TlNet5iRTIA1Jnw+urBO7jiiJuDLlWfCuF8R4lJk5M66jDQRY6p1q/rbijMHX/qYcRvk5Aq2y
CNDBXu15vIyQ3EmuPQnhqnQ72Wc6lE2TRIxSf+OKCG8j26IT57m8LMRi0UB37T6Y14EtBXVyGKxq
eMO/P6UUMeR3GHwmQq4ym44sKq5UXaAbaUc1v+RcUkX7pWHcacpuq+J5/oBEz3VXNvl2AWmQKtih
Gy7umwoKi3fWShU55WxjwtiyK6MJ7yvDEHEsLgzmvHoDxmSx4gQhaYwCQ4b3wnJ0RxnbGG0c0D7r
6L9Qx79U7Cv1p+bOx+IngqWaP62w0NPACRX9ka7qykxlpwPvr3AF6aqkjlwd6qT5LyGOB3kKTdMn
VVgNlcTLh7vqZQEqND4xig9h1eQAQOOkUXAztCmGbMSShS+Ew8pD3Ox/EDFbtaWRRcYwHdc3VlaO
fvuKiWrNx6gA95E7RKXh3lnTjY11s+kf1ov3x3gVJZjSV0dRN0io4SqCUEs6pz1Fx7g3SAPFmEgN
WzjIfMliN4H0KLQlU3w9+GoVahzExMWuTveAX1EBfNTnTZQvjR6aaUsMDJt+1YIJYIMVPAuvl6Cp
ypeUscGw2Mg1B5wXcS6xnu6m5n3k7jiBtwQOOoC6yi0zZQos2lMqWHuYQyyt1JhicB/jRkUejYbQ
hOZ4T1JWFpzakx7tDTz/VOv0BfoMJhrF0AocB47AGCJA144XGRcXBTp+AIebR3WEhgvCklT+i98+
pfYHPYJaH3QakrXt8xQEqw2LBScnwPGt7W5ab4jXf7pTIGAw7fGqmgvOntpGhFOI/J1Y0+olivBB
D7WWSp9YOdejKX5RjKLAb2KK/dUWWL1mVsZVzLudygFF9Z4ldvnjmaeMUL8Myl6KBUSHHP9m4jtH
MtUvyQpOFP/kjYZ92uLkIzRGdjfSm2KEPXYp+GQ6LTeZRIupXa6eCSygW4+POvRxUEqY3U2moKKG
EibOATVKN3T3eEcpUrE6oc8suWytoys0G0xr5JgY6g79ymfwBTEAP0ha2ncyvnogaG+5XIZSoXvF
yw6PaOouHWT0dvKIUpLRW85RTYJP6xmoKNO/d61nl7mnxG/FO83Vj4PX7frAkseaUuBG3n26iHQn
sgBAE23xW75cHXAfJ484hw+AI4OnIA1j3k8uWq9iLEJKK1PDTH16O49Xxz/noxSijhcC++dWBuaJ
hPhxqPnSpp1+NvlbPuv9lLeYoO1LQSBdUVQoJBYSrnfQb+lPMLoz50hU28ktwXt4QAdS/P2j5CO4
ZPGX1uSPw7EFL1mOUDU0UvrdBEnIzMnxpHfhq3lh0F+Rttbis9+/C0nNwmfRzO+ooRilECTffAZb
ZaBbvwc1vbH2HQfHkYJr55Q2Zsak1VzbQ9Kv7Frl+cmjl1IsbqMwzPvedlKDRFwYF0HhHYZWuyNg
3jg5vTpDi0V3uVtYrmh/zKdn2X2TzD9UEsmDbYpc4wxza3KUe0fNdAQS8kD1K7uDxPNL6jdn18KD
IFRgCazGXgCVZ1zqJdiPLod1Izo6Q+wO0ibNj/4yqjgz9iyDv0g7fBzh/mAWQvV7uOG7aKx9e/EL
+kL6BR6bpWGLc2blZjY9dQX90wf/h0mCULfV5DJFRWZJynqsRVI11F9GA/mKyLGxLBjA2gCp/CAk
z8EIw++HNf2t1QMlfwgaBSKzxs+k4NHF+jBydAR0Iq+G8eHVzc8ImWV0v4+9llRZ2zFq8xDDatZG
K8eHwOgDPJuq+7faLW8j8abz7TnjFbkc8iI6Wk+mUSpKu8P3KiAPnGYGLgsC7MkeJxEdItGjSXCI
zhjVPuR8hwtzLbJf3n31jq0rCCWU4D/lUuXgD8k3Z0eL192sRbcrTGOxXl1u8Tkd+OPsu0BwHVrI
O4xMqJsZmaEPacp5LuWuD08po1BvtbGN+jKo2Do4r8AT1aS1cLTZma9dECe1WTqpoaaYGTmJE2OW
09OR2NXIAV4QlE2QAh4EUKP1pV6OtqMGB1abucPOLHeh7g6D7TUZ4bwHknFu5jbpPt1bex7miOLm
4xEu5xejKnOVsAN29U9yqkQxGOchNG2tcNxW3Xe5Pceq5XQ8wHEEZainRsvKuPV54aqNJjqco+Le
URwuUDyvbbhOgT9joDtG+lwkcDoBbWTuw/fflVzzIXy1HvqxDyBDdE1Mlo3dXTFpQXBWVvB3DTj5
6hl8j02CmJjJp2Uwh+Rcome0q9kfj9r2mltufUui8VsTVHXNsvD7TnnzCyyNRaomcdMt0bcu4Z+v
hzWHHj0I/c0C6fVcm0mZd7MNUEXy/ghmlUjbyDVDW3cOvodiyxCydT2cNBpFHeQnqww6UKJvmNcT
SPY6++0p68EdwpKj1dMjryEr7ijo58ZZgAdyUgTRnpK5tA8J05Shq68YH6KpPZw1yrcGEemF9AZi
FYNh/9JFoNI2R47gm4+YnND8HyNJC4TYUPWbTsxvE8HZ+x3iLYUozgi5CUSlLF7saLG3c2lD21/S
Mn+vP5ZDlaM5Jl104tAHxe/ohVkQAcb6K2GVCbZxKnuUmEerElh9mGjop23PakuJhvNJtf7Ji3A+
X+Wkp76KZdnvkWI3M9xvZzt2/67Lnq6xUmYoJFtsGg3qISkpHKdO02ibOfzV7k5r/BVjrgD3w0pe
pyKKPoX60sQQODv+8kFyMCNmvv3Rt3/gDVaUnNPFYGzRYG2+H9vl2ddX91pksm4kE+ZAAlglzO9Q
jurh/NUpNdKMhJYURLOKMws9QDP4ydT3klLsupYgiPDgclI0bAVeAVMmrtEaIjOXsc+qwZs/tdxX
S4N/dw517eRHKYgXXgHjbaE8n6btQBW1N5C+fdfDDq64xU1myQGXVEuHdhE1IfHvCiEAFhjo6Vn9
kjdfCODi+Yo6c0oCdma1qq01tZElGt+MGYdwds87lm2y4vY3EmwYzW9X+z9U9JbVq6hbW081Zuvx
1Pua6wGY3TTh/Vm5X8+P4w+xArb8h6BHHWKJy5Zx7SvNgAIQ6ltohBtV1sMdDkelAY/6ccH4nOMR
WJ8yEvplJlUV+/50EJHL79wDZMcGrAw9rqywAXif9X7ypmirnlgSMG39uP4hUVZmukBnuOoowHyu
HMLN5Kr1GpGAJGUqLbXXPvlQGZeCw/kd0HH/UHoUZG9i2498HsGDThoKMca5D1pxz/i3BZmbRldA
eFJKiXYVYutRkSJeGqvHk3I0y9GbdKkHcnlXWennBr+7+9BGbCdTDQdcu7nY1xjng6vljKgVhpMt
+XRm6+uknjNOS/KnYKS3JGlkb3cfkzsKWrnUOldseVtrHdbMVecmPAho1znWzInGydygMlo2VhDO
VLsE1jkS1G4uOgb2keKuRqwqC3znJEcPJr1K0CMYKglXyTcQKfV6pl3kTrsFEcvxilyQKSwNpwOn
hCdiCthq5hkUJX3z3evUWt8uArsAWuWa2K/9Wa+jyjMQvbSVZgcz9NEYNLFByWG8TyK7AWPMRgPQ
iAdesxZdug9+0f4PeXMwVrimqNoigX+GEBy6Vlz+BJ74vrktYGqY3Pxqqof3RStosWu5KV7HRYk6
z7rsfQQMO+RIi+y/vZN83mDkvLF31g2GyBWdWD764fhzP5rzDg8pA5J3ZRtjkIIZEz11MbZWOxk1
ptN+5FCWQIyPPtgpM3gAYf9R+mLdA+M6VRGkuTcN5bjmO8IxCtLwgstOAPCYfKC7z5XttcYuR2jW
9iD7R9W1esBsHmejq+odjFqyMOcNQhPdin79dSKKyuwD1cqSlp59v1GO6Rv0nOD/17CjjIWU4Art
s9kF8WsFz4NBQ8INuplWhenN9FNwzoyS9BI25QbdAKFwMTXLTIoVkAoqruy93Dj/b+C6m7rY06jj
I6vbb7wz4jxvPvZLGnGUDAKD1WICCEwf72ZtOAaZieg0f9cNN6nzvMkp2jjxiWC9EBOY8GBnPJ2u
ZqnOotE33dQ1jjPGGb7QO0I6A+8CRc74lVr4lVhKXqzf4jymjAaiiTGiC2tUhkLXVS8JH9mjp7kT
8acJ98rolyWmsUXE2QcAEiSjTBykynAV/EbTMlfKWbITz4uMDWRWfKkoicm8nTtwuNpP9Amfrrib
kxunRNlhcdG0lOUunh1TRbPZtXN9SCSNV4ioHhLZFKr+fh0LQm2KrOfIUESBMbtm6oDIXU5Jimdw
luNo6Ohi7qs/orzuEL+xcKtS/Xwa2J0ComyqFLtPPwg6aiEtO1ArFLOaQBSmm0ta4Rmzpkjk13Es
V5Rqb+6ADzhhqkZe2mF/88xkf02vxF+KkszIkuEv1OQW7pkDjg+K5mScHZNMKSFwJ67x+a+aP0s6
Ivgwb+3O8dzLRc/R9ICRbKydf9zq2SclJDwCi2epnnnYf+C+D7LJNSqjpJXYuhT5m6zZ1gSMc9M3
tlzM44mHvOFoGyiBOhp8dgaJD2LQEgl8mfGRZdtbrdA9CZ6pNjj3q2vOjKq4Zr6n8E5PJL/9x+uP
rjq1Yje6C6XfcyahdTqkvBkj8gcHQ/lyMx/yKzHSx7Cs66EMCnWcKOcVx7XJwqhjzNDHWyywph+t
v1KEuaf1J89PfFXK4iX//47i/Z1ViUYILPvYALmOxmzSVeah4XpNn4jgiNYwhg46wSxByo6iSsQJ
6K2q28XQThgGIHjxPGCMaWFzQRzhs6qFBHcPEnFQPCbFV4YQ5nN264ECOpp4j7rtEN6NUEN44vnP
X/a6NWNPcUDiFvSPda/aqWNckA2os7ImVrFLR6gImdn8KbvP6rGqhf24hvkmgeDxmsthlN9TqLRP
nydvGr3SR2RfrqAnGQmFHkdS59Bl7hC9K1tC25cDmZt4+fIEPKwSPqtwtC2LCV37qAwipA6zXb18
Q9YnouP54cgFy/oKMWBe3+SjEkQRQqBoFDOiYzbihMc1ZB6ASU0jr3q9fEF67Cr4DrzMUV82G/1L
ujTybK/ltTcOuZ4WXwk8c+cQJTFsNstQlaP0Gblc74IwrVEc9mKSSRi7R0KZbX5svLqrnphygql2
YRufQFrDGRfeBBDltsvQTTOu6AjJ/soTI3fOFd9z/jUgQTNf6vIB0zaIKEZDH9WEq+WzdfzaHs1Y
gHGmCdaZ5IBSq1p2kXwZlFSxOIIDucfiKn7Bda7+kxROUGiNnQBvXteaeGBJgU7YBi5P6BdiIo3Y
y7vw0ijfKLGMq0XV9ULtNMdUSIPeBeW3bo9ZtIn3FKrE1B+ujertUDqtW9kWSz/7EJFlPanihyYx
Rt2469lWk2UggtN/9suQoOlVK2aqsupmp60MBPZ+ySlL+wG9WCinMzfGXyWq5s3oREfjX0aVzi1x
AjKsCZGhD74XnL9RbgbUZ/udiGU+PqXjTNpuvQI4YgUTynLIHrEGCC/jgZCnC8VIoiNWni+iR+7b
eZGTfz/MjHE5WtPFUfUk5/aYU0HNLD/p+TdI3dPTFzlYlt6d6pNjJ9dWUSKI2WM7Oj04eZVwwrpY
F2ilp3R0aXRcPB3uFGfCmI6A5KQl3l7gRjlqXqM08N3CtDAe3+9gAAJ4i65L/3go1TQt+X53VpWc
ukT1G8j4rhyTBPxYePNc4MYY4xolMOz+ek3TBR0mtYUhq0OYyBwU0S/lq3tqfCoO/xO7c+UgPWmn
ytMygmeKepjhkjb/5mvy/rx9nvJfYktQewGwa2A0xqzbr38BSiux067IMzQ7fQKLAy7qvvzhXuEV
+SevL7SpqI8Q5xuoA9b9rLY0etLrtQHJvVi8jHOSpWErsn543UvDGIZTnr5D1n4WsPCxfW8hKnf2
khKBOWQ3rwqvoTlRB1oye0cQobTZpZ3sF48PADs26+RgrWJu2aXqUlVVfnb4IuzS2UBOjbA5TzbY
T4yo1GyzGX3U2RlSt64t18i1ZBbXA1+hi0ybalM/9H85N7AFQVHvMg5ET0yAQX+pI5SBZvckV82u
CodzvVg7jUqJx49jegwEE79/+0uyUIDtUCD6dncSzDUeSqeRcTy5ycIcILW8ghQWflyRNtvWaJKL
7LEEEQzWoxgwagwSfTcxg1uKSHThc586bGC6LckSvfAm2qMK7c2PwisYJcXVDbgjXGJheHGg0wZ7
kwKnL5QkwZ/PGM9+LpjjdZPBaRV0wkaTgST2NFCuElvzQLhvccv0E3IfhmzPfNNWN86jNnLnulwb
if2sqQpVRtOWP6advs+HYOz8juKhPmpl1rJnMDC3qupFcdNbnPlWd/vQlsUrSs2cyfCzzlL/zewu
1yBIcCfmpNJ+clmi3vmK1cjo9+4EU0HB19mRN0AtVxmEvLDZhRyZlG09gC/KFIWF5r9MYuepm31c
vN8lPfG6XsSpDGjbcfU7Bg4cybqueksevxAQxDpAAOyJqgMur5K5UlIxCienAmTfl3FCvUyjzsJO
X+gRmhadP/S1JtDhg1xrYcA0yPg9vi7Jo9f6LOpf3Ek3XZvoCiNq+z20DClbC6bOu1WGXyJOD9cx
9pjc9TR4z7UDIplfuJ4f17J/UmvSCZaI1SYlkj8ZN7qp9OhLoQu0qDTDsVYsRRDtDoOvufl2IEhF
iQLf1k67ZYg+EXC0DCW3C4pXea97dha1V2RFmPqDYNEJPuU64YDP6lGzKs6bx06YNpN/0h0g6aIc
XIe7M9aMNqeTX0xkQ+xllfxaBA5qJcf5yLPLv0Y5yMaMibfFKVCAKvpLkmZK/RYOQJR2GVl5QXxk
v1gZlq8chy2nzqVANp52ArvhtI24ntHR3jhn+QfbChIpBVQO43nX7hyNTeB1VP7vDIhx1U8e8kO4
HGwYhCMq7j1/8w7TD7HbDMepJzzsujf3VG9W9OFOGl6v/yZzGTshVcafefhGfVYwRoTnS2GHPpjN
7C8DRxGYuLeJYNeEXfG7I2ZpuOfv5r+n50iwSL1MbTlB/nt21OT2s5qJNWRSELY6lYIdH050cm5J
5gMqndav7s9gPJPzQVGdvmTp7UJycCpmuOqhVxVIffbPsCPqc9mkQRsEue0qDFfWcZJWvaUCReBt
LxQfEuHE4pJvf04MWZSiwNVn8n7yBpoz03Xik6zC0TDnYJru0DlxlZLBq4ao9omfEUMNQWWjkNRj
A889WArKKzxJZk4/soyBNpVj7fJEKWoGMbn8tT4YpFMQN1Ace8g2WTE9NZ8LXvwop9/usk9Fiwc2
BqTzUVzgkcvMKtr2r+ebda6gaOFRXikvu1xdkpHvncqiVLqOci7/xLypB491HJI4wosKitSY6T2C
ZOdWCjazSsehdxVGn9S1fNAH9xpDGRpxOrRvByfk26xFZbm2rfu/xBanhtTXv9fib0jtcX2LE4lb
G9CdvfiRkiFXgbbSmkxOF9V5/WaRG+Uhh3ZKjsIfJ536uAEn/PrrN1itapfp8vpwvjwGgX+d+use
qxZBkE+vBDGAqLR5NHBXS3Neg1zoEoh6cIDLJ1DwzWAkXGDaJv7ltJ6gcOXsWnShESc8+pvDLc/P
MGau2HqWWwzAitIqQlJulXETBczlhJC2skfBcOnmb7dvxpd6XeOGCczKrySOak0sP1BpZuJlykyi
NbDo7VxCigS7oRsPoxvRFpvUCUE37jnuQZQGPspqeRQCQR4+PbMu+LTT3LIXKClQPTtDnrXT8ua6
CCfLcNNqsrHVg9M18cn0mrTo99jY7pNiOt1R4/1VtPky0go21hKFdVnlBzaLyj/naNvWk8DIpOLh
dbR4NJY4r+IxnMkj/z323t2uF0lPY2QHNbWlBaAfbDB045zoieF9zHBG+LB1nFmufU32/wCk2tjO
1RkJYb5BDry2VYub6nkL5Cc/uB4KUixe51gZMmovIPBH4didjQtVKHCPhcGUqFJ6dKylxUCPSmMH
TIAIKt9pV+3KyXBXjbpbZ5EMa+htIFxQdUMP7NtL75KlAH4o9HWk5Dm4o936peAtx+IYyj11nWk0
TwNDhDFiwtultLrFft7+A0ygnTJmmcjjg9D3qxZRYyYo/CuA2XBgGrUzPmU3ghJZoBcZs/fUpTBO
1lkI5kbxSyNgXuTKTJRei4rkNWAQ9fFfS6Kg+DkyJfX6h04spRZNmecCPMuiJ4Mh3GL9DoN/JAmT
6nAtqhl+TSLCyurge0NkVYXCJWxBIe701E63opvsQdyqmyBk4cgQvO7rrnsh9RDGmnEdcAXImNR2
oCm4FrXpARkDuIjnXCskUbZAXeCEzPKPJ4eHXc+EG4ZvBkhPdoNc3mxUoG5kgkDs435Munr0ZhyW
n1eqrpJm/tVjDijiW87TabVadimL9eWv0qAOuz1UYP7yNYrFdTBZ8GCloIZRvILDeeT72fNevQ+W
KwhFCNxC3ZwrWPQkb/cMT6mwesGKWZDKA9R1XTM5TET/QkxM2kO6rGWe8eha7W2MF0Rfsaz1mk1y
7Bj4FU2PqjpGxamL9g/ogfUDKZ7691435e1emVlhORMSAKxWpAh1egRGM2u4PaAfjgZi/LbWjoA0
y47+0kP5dF7fxVmZUDW7Zrba6PFSHqV5HcYZoFlZfgeeeeWf4pKWrkjIGTFdHH3qFsYV//R7SAo3
/bEXgxf83zb0+bOaH1ACAzoi51wVYORJHoVm1Pm60tzDnh/H7XWdTU2J1EoIsBww0WOcikmNYspO
B8xh9Ape1/sBDYhBkIy7WJmfwqa0rXiNQISxVzLXX39y5oIqO5ZEADOBeaX4PWgyc/k9Sm/VggYx
UU/jV3gyuvWBkz6GCwsPXfUZCUzAkdungVuG96fv9k07CuPaAYoM6J5Fd41fHTU/HU2WGlw8c6a4
EzdbdpmyzGZTw8VqST542MhIokrltUgC8oUz9UaQbQ1wC3u0t7wLGHkCoAPjiCwXlYaHj797oVHl
Y4lHnT94QnN8do09ughLaS6PT5RdfU+y7SRMkX2KjZo9Ml5ZYhUPiYIwRIoQ7FOQpttEF2HfwES3
jnyBmteAFsONIz1uvldJatX1rhBU/uxywvnQhNoc2En3KUsLmt7alDBMH1TrHrxWvaVlqmTLghFX
SGU5QulPg68lJacZmtYCnoFtr0irURlMWnsWqTw57EKsIqr3AEavmOFUZAExwus3BU+TQRJrRDnC
ncDjsGVGqax32Bm+1IEa6idwprgEAz3fO1hi69i+T4Fhuvf8OaC7YQEKX6U7YdTA3LwBk9djhneV
FlfAnBiJJv+1X03oxn+qD0Z7vpx3g5whN+kfDbu6FCPGUjCv+SziAEb2ubGm43eQZkwyiGaDge9j
mNJI0AfxAI/LgAz+Lv0O6tfEyUs7pCAEWESGmV1LWf6cUuHPzzkL4CsB8Aho5i/ATaxRA5AW8e7p
ktjjwjUFut9P0wIevi5lLlDWnOdiiqh9XZLaNnKSrz+UH+tOs0e9O+rClHeqItJqL8ahhKEUhhAh
1XTiMFyjmsnLK4P/x49IRwCQBILLqHRbpTzGl7A4VyJo1yG/ZbTGc0a5poVFp463kh0cmfc9wYKc
r+XWacfiVznPnbM81jiQ0KSS6LD7QmJJVhCrcmi+Ma4ur4LtmdA6/6+tQ/FlvFDPEfXxDFhRtNe5
L5pdhsrqe4MysciaAbmvkJHBDykaYHU9OkVyM5EGND3llYKoQpV8v890OfVTtxrRPoWQ2k/lsW54
zn7SwXAnBV9qOddnLvZgq+I/nBJ7ubjaO2DHODb486uVum1Ih42PYPBR5+UMtSfoTi4aNvMwOHh9
arf6RAJCSIJVKQuLZAu8//L/tFfRf3gdb+C1VjWeOn7Z/YOFs6RKomJwPGjDvdlbLFPHDeHGhs8v
GcrcTBm0VY0M5YZQgbL+QSNc+NCQkEB+jZLqriutEX1hERkLXvrDCXY+XrS3kawiaQrzluWfc9iC
Ai1jWji8UMB6TTHOPcye5dZ+MZfzJlakV7RPdznJPvB8CBHDjbbjRmRXh8P0Rbve0BKVajO8BL63
RlT9VL6c8YkIbk7oxwiD4yhV30AWJ5mMaQTCG9GwNv55CuFLIJeaDGcNaVk76lSOT8mievyKoFJP
lq+z6Y/FtIBAoKUcEPOMhQqEVq9fik6ZySRfKp863d5heaLxU1vfcNpOIKlWoXO1IlfDN2g47nzX
I3LFk2CFu+W8z/eNq4tuaY4vC/E6SaE4xk79MGmcoNgPasezmO+BlM4IRS6NX7E8pQVyn0m9HVxk
NYLxjRfo7BE5gwotukykvYY7fBtvgl3WFCWPxuFxDtyY4AeAa2q++zKGkGxGZiTvPcBp7i3sJder
3mb7X3EjmBVEV4lV1uAvsYsijnifo+nmjLljZmQAI/TRTMQgWKcJ5quH8gsUV8wc8tfivX6xQQTh
5jp1ykWtRsx12AR3nb2E3+Wr/sEbmfK1o7khJ94CoFQcRsnRkLmVeYElRpADxeEIJCAW1QiOIXbz
6leUtY52tZ+DontVqoscWbAPmywgtBsJ82J8G04ZgOhTNtlP58pLAP3/gJP8psMKnEXSg/RaAlIF
8BgmRaMtHU4m957YTpEv/xFwcIWt2KKZw9vLldMUs3gqr4lMuhvrzv0AHb9QKB2Yg2JxzhP15GIE
TxONUwRSxnmJSJk167pEIJ1+BIX1ktvXphpcVVygNe58EfMsUonV3rkg0x75CbTK0NqhFDhxPeWN
VS00JJyZ3NzaNtQsyoJ2tgeiJjmMyQTnoH0MnfkE/LxZnNY2fHKqIEbQidjzynxGugdqm8OAHtZT
redutLH0/AwjVr7I6Xp0OJk6tFlVzaKMXDd5AtUABymdo/LS8fknEekj3NIIjmGftgdXWS4cJVBO
bH/u/LlR/d5xRs5zEl5K9amPdUNUgW2X5z7ufo6+sD4wwC1//SasDpqFW8zbTxUq4dwaxFisVfR+
sU21JayHOhlqXNgO1FZT0C9ylBC9/qDcspB8HKWAUb0nAG9e7JdLFbsCLlPnW7lKugbGI3m7f1fh
v9X9mSxjAesRtil5AC3JjP5SouPIKPI/K4uGBq0OAemDvUXjIeB4knzj3kzH5sLbjG22Pm4FVfda
RXiqvNhKnf8aSamEeS+63lxehFSOtNiOhNJeF6c9/NPJ2wjckcveEYahqfXH36AKmcQmGkTQLTrm
9mIXMKve7I4rq5Bb96wWq6IGJh6v4cDW9lQvNTEN7eYZJO/DXpn1FG9XCCyB+A3bX7jZeT2Ux8qR
QX6/b3Uq5qN+j6aNwfDNTVEOszHY7N9+3IvVm90nAWI6DlTE98ddK8eeXJh6rMAoyosJCsVMCDlM
yRSdnsumFONfViam5XOffFo6noX/gXsLZ7Rqwe9kCywZMGX4sH7stgSJH8FgWjEcyIgCmlirgqAy
7fA5dzUhorHZaq6g76t8GkjM6YIO6r8ixwWb3aJHKT/luACMuMK4LiEw98uuQ7VP4ozT8lO3AQyr
j8qRSAjsDpJqeubmhu1q/GBRM1G1sadTJgLBjrQtJS1eDK9zXcCi7z7FvJZkCiQvOnST/zLSpPuY
HfDkw0dF5qLe3+213niGs3ebK7SzwIH1ITCqZmRdAkB292u1AMMgB0ccYiv9TwMZKnfVpKM/aERd
DkiDWXx+H7o5vWW65iqc84xe2B8jaAg7aKsZEZsBtAo4U4OlmSp9XUZ++GvlPlVIjr7qXlU0K3aE
zkFP0oFW1yUDHvxyp7sDXqAi1QnCFk95AgLLadslbBEO1JGG7EcppK1qiAa0UWN3YtGqpgaDqrjl
XNb+7FFeeJcID7VXPl+rFcKk5kEXHCkEkNEEp9tUaZ42Pr/13IYW322O2fAGj7Rq+hIvs+qLEHwW
RXbJBbSFOPkSEPZHG1DNcnOiGG698qTz/HOx/UnLeyaBwPmwT3gYUiYMdBX9U4RJNaw92VqMYhe0
XI/YPjWe0Hxwfka9mOaop4dBqI5dyBgn9jgcLfp3oV4hrKMl3u230FaL9QZyqwBdkVZ/1R3jvgEz
bSmhXXgU3wE/NO5DFBhQXN5Ndz9+cR67gHr8OfU+Euu/cTIi3tQf5lXR+ukG+FBQr0PaihjL77Ut
/jTBnvqjA5LgZEWQjN7D4VjuFUbgYQ0psDcen+44PMa6SSDi4ibBTHAi4Jte1yiP9VHEI7DOoHJR
DOVlydbER97Whz6N+uPBkt8pB1sGpYfpjLz/JXGHf1XpXShRJg7/PIN7BEIkMA1sojvKPiBhxAJu
/s7AChW+2hqQ6h024+7dBmotqPYeQt4hLSlDvp/T9RvKmt89j4fCMBGApTGsnZbfhD+GJ+s+E1uR
8or+eqzdVYGlX4KuNkuWFicmU4OAFtNtGQklakVvU93twaeygYWO+D6mhd9i53tWFUNBABzQ2cQQ
3j0HGr1Kry092Cctjit1awm6IyFzs9kKfllj3NJeF4yHe1JfI/6C/xRVG96jiwWMYVB8HypeolzO
SMCNesPFG75nbOqPvnhAZFJ9nRuB8GXHR2dSKABByqiDmCfjCa9BXvWju6/8mSJZZO55iO0L6GNe
/Mueu6zgJ9BEDWIn0qToVqmIbluHeB12T73vzCGWrJhfC+EUhiFhSq9U29ZWJBN7Q/ISAf1X7qq4
cKpggLfBqcMfGhP3dS4o5w8Ov969/DxEX7qxwBm3GavPu5KsRLSzzW1yeaLQL+hdTzO/CCXFFUGl
s3k5E+3eQZ5veH96ujh6k67Ao79sWt7apmcxWOlslAcEccGGln3BSVEjEa4FMow6vaQWzJqisU8I
hDWHHSudK5x5ydKan8m3vWSpFtB6Ywbf1J1s8ulwIybXm2jCgdEkfp+8DG57Hv/eEyJpRwjpXkgH
oPXQWJiQUflgeUHQExltl2ZWqyG7JN0KrwVs7hCqdHSaIzM+OTTxkeif6pUNBe1z/RY6Kf0JaNtv
FKErGzH878PPXO6eFqAy3PXRI3I22q/JSTtBcjLTPfJ4uAaU2/NJsqT0NSIrKe8uEgPPB+X7VW7E
1yraTVKjQ5c0ttWdhgJk1AcIq2iH339tC4+2O43bdQ1cDRbd+RQOanLwyMmTwQmHLXApeLf4lJ9S
NzG/z5VkAROjVarl93779sfuNcnON3BEs4Dllz4clMeS3pboDuA0vFWGV1H9DR+bQ27wnomH7sbB
c9+rMeNhi3cbtz+HtqiHuRJQpaS+tDyN+fGhMWnA9iguEDEd036BJ960TYZQv5tZSK4P5o2sbq/s
Azus+PBtv85yvS/QgLvzxoCPgibKGUJLaHIeRckQQG4xlWG5p2ecj75ydjYxbukDk+WpFhW1E0WE
muzehcxwmFCQ/D2Ye17l1pFlP82z0aMboQOWvyW8FDTkjdKLQNYaHsIzazlRxc7YLRQfzpH+51MG
5iLj6Mky79jSBQKG2bB1Zz1K8ufwl4iImWgfT7eYd5FuK5mnTEAgXszNnURrB2HzB3Xath0fJ1IK
uztL4bM+FfXHcDAkFp1FbKyEQ+LukotE7gPrJnGzIaPRsLUiIr3mGPQayx/W+GAs9Qz8QVKzBVOX
iaxmdcLTlAFJVUk7PqIqMy5iMAKmmBoCTWcyM2uQ7Nk+8hkZ+JYnW0jNBRnikjAf5kGjPjJd9YKC
9tu0TEk0Yk5n0fnoe6LaXgrzKijOOIdfOjUZ8pmXLLBNNKjBOTj6BDzWN0plXeWEu5hb0kNf18Rn
QoWHB24mCI9a6J4/5W0CZVjy6eZwbNzKsYm0nDcL88yjmipx38nhxJHecY4Pc8BV+rMx8VN1oBpy
WdhxkQnUeeFZDvg2CbWihyMz+Ji719AYvO5wyyQO/sjPkU1sRf6O050ZiUmt8Xs+gI4ecWa8WSzc
ddvYvVkl+okt4KjJn4siisL4DfIN2edYx5dkGeNwe2gDvkwRXyWiOmMLbHD01KjPm/wg8N0Hy2cg
HPvJ5VCREfRS0OYTWbs1oKEeYwdwQhTcPgupJyXRHrPdBHsg6crIkFpCjhvcSzCdJGRLgOHYNufc
s0XgImJs81eHtO+AtdgGObAymvAm5WDAoKrCVUe050gVNKpFMzO8U/0EdvbAbJniBXnl84v/Tdoh
h8uaCgbAhD5tE3n8CfvLKkSDN34ZPX59G9WS6D1bTjKN9arvWA/RJgVmZMqsVFwBq8PXWkr8OuvC
u+1j0qq/rIr/6fsV+aPNZ5TvyQnFF8o0gptH9V9AFGzD52XZpGhoGh3bPg63F/hyYtlXXP0C8M3p
W9+BLDpe/Uhas7dirAWfDx1VUIAMj3+KMlCBruUEa7ONQk0hUHmUTmeURrRkUB+TE73oOp8xM+Nf
TnlQnr+eRCaXF82OUHst4wnPwvhiC0tORCVhZtxCbiA5d8te9+MRK2eK66Myy482MxpDXQ6VD/6L
PdUuY+YAzWrpQo0QOen/r9D9uvjF/s9m+ra++cLx3bmMrCCMzXlHlBhpPQpvpVFvYNF6rs7ufT4l
ms2gTzYJsjtCr1ENYLm5gZLt8uluDt64TfoeVDy+1rCktxOSkLD53nixXa6NaaYKomY9bxFr1MWQ
FWcXWDjgQhc/ghvXZ55ovKiaR5AaNR/rqIjC8d079TGdKnQ3qjYNXpuCcaFVolvProswr+Q5Vzrw
gW3tgziEd6Xb/NZ+HVL6IxZu2XU+Fy96+3jSLdPm8FqtUPMqUSozQUDn5wUeWpz91YbkhHLhUZsV
TW1aLnxTCXZnsp5JvR6BmwVWOpZnc9UAGxYl58Q3e+ESHh4n41/8DXiwQo99R4ispISgPGKJHkqy
2P6nDwGKNUO8ET5/W+9L5qNhAFw9YM2li92nY3UuombsB3Lo8KOcNwIvrlqHwfSeKIgd3EoBYTii
ktoJe2Uz7h182SADTj3kjHWdf8pNcUYkNCz4pM/mVBKMVc4BK7LmY9jmHwytsFxXmclLMTXKcZ3d
YT/VmsSbpiLtU6E6Alb9ziyJ5BvBeIMJyfcJQdIgOt8fyvGFa7vSJ+TzZ1mboXJfE6CjjXrbWkFK
GUzHH/fTIP68WXyO8+r9OqAgXsLQc0iU2/x4EK3Is7jZjJMd4XwEZfZpwKwvf74WUsA0F2gThsOk
aS4LBYhy513+PVZVsFTyaLtoDFkn5n8wWnoDCKkNmBvZiE7t0s+5HF8+Fi+ghusCYRx/NmR34EBf
ePi9Aq5ps14fU2WZsPEI1yNsTSJxnIqPv2hUhuhxiHZ44169PfoOTf8zZw1HpkP+9eHd8kODPt6I
L4MiqYrIKU3FXx3e7ttv5h7jPcpzUZue/AH12k8iOHipbnq/l6r9hlK3jF0Xq6YtksqU//oswIEG
w3gJUnQjynugQdvptRcLson7O+X7G9Vu2bWoN6zo0esDiBJPPDOXXlXyrEuCmhXUr0tdUNUd2CT+
chTDA6yt4k3YutNyeTZZCz3vMCa2CSWuCHMPibQWSC785BEaxWkvM+5FS7dG9YrFRqV9Tb60Cu41
SeJzVk7Hnywm9opEt11VvCxxoNeb+ogVAbvKFkL7VH9Ib1PxecgpD70YIgC4O1iYcbU+RiApMnTz
74s2oCk2A1+9ohO0xMbwyf/vvxOmtgaTSLeSFE98hGp1Y/aMphD9iGWTr1kNUhqRZvkcLVmn9TbS
Q344BOxsxP6dw8098hC6cKtA/CVAYxG638h+L5J8RVlLl31IdsT5DqHSbjgdaLo4ye1omGt8l0F6
AQTGZLUAesJfrwCohSFJ5EM3NSPlQA1g0IkTJ8HgxKu/ADL9iwsH2V/8XzCxgNPgNhEtcmlSukU9
ILisU5fOxckRe/g4QOVPzbWaD6D2ZR52EKgUi/hht7mRKdgBf2/AucpKg3p5tVTqapJ44UCGIBOT
4E6rY/nUH0MVt7efeVAhS684j4edDabXGO6aRvUALl4/BlQStEEjupmKwMOYXvUMii5OigE40QxG
4y/XtX/zEpwvQJ5Z2PR+Dtbh0y5CnZTEBRdaD+8xeG8yhBxIrpwZj87H2XOsO9/iIWU9iB7dswbg
KiA0s1fExDAjv+JqdBkWB4ydrcDwXYPAkapY3Qx3NhbdxIPSfDo2LaO4j1Pz/YDpBPc/dGRlqpHO
DREmAIyOEgPBaTnTkrK/8D+893BLDxg9W5gTtyOiyoviZ7H4OA2En66Rwl88+za2A0HxNfbzhSjP
CQGCqwNn8y8zOxAW8i0jYfn3JCl7iQXKgJoVjsOqguQLsGFlx6tXZVOdtKYrLmn7bqy2C4mau3Qh
gDmMD99Q4RQqxOU2auqa1lCEtjLvaFg+EcEOPtaFAcCZC8/t1TxSwuF9luz82wdXeA/a9GSUj843
DJyQXott8BqaiNf8xZCKolWhixnux+OTss4E6s+yrqs354QnxFrSumG2rTQv6+qJ5ILgPQeqEl6d
ZzWyGnzDqwLEOPigRusWPgRBUnKMMBlmUr7ucwz9v6ZBT42zhyeKBYFQZpVZMFAptHffE6TG8XaN
C3OgoyHyi+9ar8kI1CPPHSm24+rnoD24aAcjHfDinzP6hwp3JLyIKf4divEtVLriXQwtQQRmXRnY
XTl/RLTgQtbj2GtffoTZRUxzJ/sEHhVi0odcfDypYR/Xpm2F1K4le5LDDMc8KT4DmQiX2v0B8JW6
rV6spVkI4MII3PdDKkWpjzmjULD9csZUhA7NWwoxL3Ix7Yywe4U+YYJniPaIPW7tCiReiyE/hQ8y
a4F0Dc1fyXQe63IvkhXdmuCITYrs34c85vhQYMDXmQ4r/Yx133SIHwrhRv5GdGhgpfZqCQtiR/9p
Lew8UqJUJadQbRCLWdWAJdqwgr1tXbnwKV0ApYUu8wugw4D/lbeUYLjxlkqtTymLovPW6/Qx5VDs
F30/7ohD056l8AoBP/DxVS0JZBIRsrB0wFt15SBkir++lLH6pQvqZ/0GRzMzV6NvWAjTm95CWtgV
AngWTlkmPluO8DKHBwySn3i0yra++j/YiSAbFPGxBsl8b1YCvjFH9/b56MU8ZJVm8HnpdenqCfZO
4+qt+pJfyzCtfTS75i7ODs0IpV5+1Y+982zof3bLUKp/7TLrIjGwmedcg6zXuK+w0FmZhYgNnte4
JWmKL/TNb1OC3oATlsIZE5AkUUgg/pdraaMmxUvSq9FOmCVRTEUyBj/7ddJvIVfsU6DpAhKmPVAW
gk8esELkclS9ai0OYwpe53qzgcJSJFQIt3SZI8BuN/ma5gnn/cP0rAJtUSoR3vnBGzvzR4LX/om6
blCTWbc+8IrR0sLAf+yrpcC3YrU3HZfs0DiNai+66oF+iJ4cP9Dj9FeV/6ZhFuNaKmjavTexsLRd
TQ14TFBqFCI133PeCM0LVaZ14UwvYiGWVKIHP+k7JITZg95GI9JNvM5RBosv4fdmlOn2SB8aPgTs
QKvMYtLmLeqxgZ7LM3jhEby4xYdcvsqCnPY6KKyVMMY3+QTorDBSqzhngxXoSm1s2J8TS/0lx1to
21/8BcbjVRGf2nx0BcjreYvDF5/FbSf4BWuutKVwAzsy67CrGPkBkYT9tTJX/BQ452pQIrX5D9pk
VCnDplD7gvT96fQykRbSvGH7iI1wqKu0soULtFkqwNsHGEUfp1eFkFsJJdZXIRL1rlEMQy94QC0P
27W4yF7mbM1WTC4tGqLDcZUFmwnjcXUqk32t9nC+UvUz66o5Hx7OQ6Qba+WtDW01SBxdQkhfgjoE
GSubIGQg2TP7cbjF4rb5hDtaoCqvaoVH4vVmxVAf8wP2WuOOtt7fvqXqFu1aDiEShx5z+Xld7woT
6oiF/OwV4pigjQ++Hkgnr86Ms57ZiXGpP9CdWtuLV+D1bfj9XbGV1mCPXe6l7tyI/eFyVRquqkft
ntqQtFIvkzRTc+ngRw63LdK2oUXcKN9WZkg8rnbiRBjoeNczBbBtDan8siUwSiwCrtN0PWwOlN5N
8VgfTyaK0m4ykZHj5w47cK3yscJs72tMPGLVfrlB32y4BCyfU/ZDoP6ftjg021/nv31ZSPnl+xqy
DrK3vh2W3CMtakLuG1Mes2iKMVS3rbGccAPHDfsrD5jFxr3VsrKpz6KdKXsZHQqjjW4iY2DILtnS
iNyejfQvabfQR69+wwtGbRYyyhSTWaXuWIdEC7bcYNnLD5P9aQ3jaVRNzChbZ8UppQ+FLvH/YE3D
LXGqja/WF5IJCzeawX/JLyUd7qr/pxont17D4Dc4IXLY1Na9zxjz/aWfpB3afDRHLvPQjNGehey8
iXX1hCuX/sQKI8QBc24oy1a5xA3pvCV7oSj4cx6zUeDMLP8Z3rqJhz0Y7fly4+1WcOG+M7XXytsI
hRAfK2pQ4khxEM4nBpmOBGyYoEtrZQkCmSB2Rqc/U0U3RRwCoTIBsV+BKqh+H0yp+OEeMtnxspGk
eL8pmYXAKBJdZHYk3n+pY4Xb//+QqtzhshIFJ7KNWiy6dKGPHBfNrrmGuLfyU9qE7kqhPzQnh0FK
QZMweqmMXpdArbvPZe9IuQYoV853ZlikTdC3HiRfymY0UmB6cSvzwn4rQ4YEhbocuxYptsg+F5TM
+88Nzep1wRLwrhPtO2oxb6Qu6M0M627cx4SBZ6Jt7yVyjHfhnmMhE6Rscv0dhQCZLISZklEf4uZY
uA+rtqlu4BaoUMnFnFnyGCypDkpGYxLSd3LrExQ0WGNCgsWpIEca1sNDOZsSWVrm0ax4i2rReAzp
ScS4ASZKL4aNqmn8av4/SUPP3CAZI4P5i82Dp9sf+/IjRKJfS9wt6e9vdJVHd/+OGqPFGzP+OtSJ
JiEeOLefrzcBPMz0tw+JY2PkSUNN2gdPoBQo7kah+49deplqjUUvfiey/predwGOFuJuuHnmtWmY
piG8q04Q+QlMTgK4LKIpYgvh+WHIaTTeqaUMnfP7W5BBweoueG4P+pa14V/hx91L3PYyJ1tIePei
RvPlX4Xhg+WX0VT1ww0OPeqDhSV12jp5ah+Ntek3x+BkeHm66wpVAvGRhZi3t/7duJgw53YPfpON
EOG0w0ltuh+qYobOgehCUED4126ybc9qWbG7pXXavppEWKniAL2qhU/yDfXSvjftqjKb8tz+tztf
oddm1X5Z82jHKwNPMpUWUDEIHycbDYBJDA9j80ZI4oDbuEC21Lt/TLCr/exJyohLwgJ0nYYgPu/x
Q96K4H+2mpifhwLcmtbEyNE/gznPLM1KpoW3jNMqFP8Q2rzsMtoQ6fhyvuJEZLT6Y9tQnQVcvhK2
eVBz1rwn0+kP+1jJ1iqYgy8J1iLbApn6FqEq693NR1ij3eUmUvEvsniBYiNs+jyEGYeEdih1ViK/
xhkAHVJcbVnBlD3Xndh8RxKyVCQyRjP57oSF3Rj17Mx8PZUYHUDKtLmLELLNNnuVyXc3B7kyDM7o
2aTqkxyMFEV1TLmown6W3N0Q+TlaupxBwTomoK8jjC4Vmn85wkfAPMaK8NmU12zQ0hLnReJ+zJ/Q
oDQAVAWvWOiALj5AgRhWwcAfx+ZT599JVL6WtSrvwrMfo2VoRRxMNb3N6ziBkmL7M2ftjLi/jTZL
B6Hxf75NDZVjW/3CaEgUE7nFoIcLLg7AnviiIVKjFEUUopqSAw6K+lQv3i4taYCGfnJt+5xbJXH1
mX+Q7m3KzTqbCMAkoLOVlqru4u8Gwot5lrjwRpXdpOjzTzm69lB+ijedN6jJRevTYkVAAQMjCCnS
EPgYrE4N7JvK/0oV8XisWaBylsTHMjK7wv5++iGAMVtTuUJhXUt7S91gD45wee2hMHb7WZW9Spew
qGBunILVn7gu6iChmrkvK4/BzM2QKMxW4cOVls/1LLoPkxbxwiSUJfSt/K7lTjLRUxIi6yee+Czf
hN2HVMCDsSd56mzzHo8rbhvplgprjkD/OCIZuWwx0cQsBCH3cWU/pba+4SksIW3YWXaBkkRkUGNf
OeqerZyo/KnD3NMaIRqaWziFSuOvSMRKwjpPqWVNwDkA8iAsoEGAI4LBhf0liNmPTPq+dVAbwlZB
DRPrLDaxZS8RX0gGC2FtX1jwNmC1buFqc4yT23H06faNvpnVvGXxyDD5aA+Q5BSNmQQOD6cPCa8T
Ee6652Z8r5ldjgsqcE61G8zDn93AOLDpMuieIXZfaWiQrGrnDxDjmY2ubY6u0isrh9ncP+biQtIZ
7NC4rQPjtgkYMaBh/jQ5/0rPfQRCBAexHsh19rZ5cK1wYKrGaaxwbist0UBGMtKSh7dlue/Tnotz
9NRwD8Rfo5Xi2jQzOQjxiPCb2f9BNVAY5L6cdNHgjr4nzGq+LWFnmki7IwoykBdttdP9kC2Gi5Jc
bXC+7SeMw1kAifiwHy0l/sDBrH1rkyT19FvCSIZD52anWXgCQfMue4HdRDmadkg3sseXL6aitHFf
2eKhqNuXvsVE30qErj00luR7kUYF1juYI6KE6arhd6LFbN5hHLfW8sy1clir2RHbquAGXMJj53/G
TYddPoNeAcpNON4Ey56BB+Hm3SwPmgy54KIE1EsmHHHOBi2W8o7/Hpx0SgZvVU8cuLEpTNL3yq8U
WLpAlfI7S4BkQPKGzNuc21oj1BSYbKM/tiQnLiVE0nwWsSmYbx89YFXEPt4eoZ459iEm5vVYt2hn
CSFpJ0rRM/7jQV/2dXyCNxWEjOmmIt9DRhETNkOvGga395O1RSNDWP9vNqQDFVDxUCkKgZ6Mf+uZ
2vrJzLEFZ4QtjBkgbhHrZ8ltL8ia34E3KUCA0WvZfnwe1Wk+neVb30i12HYl54uLZXGL+pmsJlAy
gBhvIukW6eDOaGQM68o6koZpOpHMTCZm8cDPtJxbENboWsNngDUc3mGf6J6/FKyWQ30hCBDuECHl
XuIBqDw9QRDEaSWHCDladQkJf7wSQQD7Afxa+7l0NpfZgcK7Zr0vVcQt00BFMkaHRAiZXgrOGWF1
rQ1nFEtLRu8IoHxy6N7nUQUcwBcu4ydkIZ9GdHDMNkNoAtHon9TYE2CMh6VImDLbnsYq1oeFFyJ+
Xb7R4bVdo/IMQnLUnMCflKTqpI8UmtWwlecTPXtG7B9g9YBH8dAFmF8qbPpnTPcHBW406/X7trZr
Y4cr+imjn/4M482aEP51u6Y2hVcz4jO8QwBwFq0Mjo1+leL/yZD3/wtLRTXE7zRFiLF8aaDjZzas
BEOk/GIGZ0XQ6zxKMcAlFWjDKtNYkJDoE8CwBtL6BInIKD98n3aicd6DURfhNF20M4UUXi1Db1qT
tUQ5esCva1+i96BBtnLlJvqaY/kVGTJi/yiMddOITu5A4jYp0jpoBa7AfnFeAdRRIdqLRi6nas69
BNe3r16eJAiDuLdC/pMn9IW3HYyIitugkxFHZ8C3qqqPmwkYVm32xVC0/dVzCqu6uGum5ijm+AEu
00QVawfEcI/Bj9uWv93vfAz7y2xe6cv71MycgFK819Qx/uFNQ1UsEBTdjM02ZO4kP2FJK2glE3Gs
QxxyfnfK3dNybuQKsSHCTUyFryq37891lSRwpErfmhQ/MmSSg5CV/HLociN2OWfcTgZWFAQZNuUg
WieXyetpBV3P1jTSsHRi6skm5YlBL2E5yIWVbRvrdknWk6qy1MthuuIKpJ6GUPdO45tiFGbvzm/l
q+LGIFxRqcGadz5SoHHYD1pNHr6rGINSGs4y5lZuyOh0H6spnL1o/KvHzzb0uxkngDuja7y7W49b
2dIp5SudlHdFY4IA2LXfpY/2W7ZC+BUlf2S0o5k523euAODnxm1TjGxLmVsaPpp8eg5a568+VGMK
CrHzaDAZJ6KtezSwwzEo0oq5aRXfdiT9KeVJ6+yGd+UxPVcBVN3qhq4jE8kmoCmStVhpM9jfslrK
W7H9dEWk7exrwMNKeWWTO0u53crSO1xPtCKAsI4UP+S7fXP5SLj1yy2hNZElsl51mtf/EiG41Eru
JEbrPVzRD9hDmATQ6+ZcbNinNq4EiycBzeZw84S1eOT1tXtOQSOvm5FywRG+UHT7okFae6DP5Jtw
fktFXn4EOHEOSpqY+dnaYDjBIdu3JVNQlm9M8/UHxuExcMKgqz2dx5qbHnoLi8VM9fs7EWCFqqmT
VxdOM2mQRxuFrzrpCwJsiMJnabY1MCI+6WIDlNnwABcDfLogtjd9QuRIaOj2toVrYsB5C0SpPNZf
klsKiPPmZriKgw2RnhHy02qRA+dBoJJ6xDFR1cUsSX57r8tmeehhkvdf8WWuNiX4lN38sca9vI6Y
Hgvqcgm4NjeNTfZcbesjGMAXvLVSvsB08yibpvje+xq9os9ch3DtFJ2jb3FqVBAAT03VNVjHkufr
eFHwPFwaBBHOhbKSVAvCsnetJv3Et0rTbSDKzJ0TMZC9ZGLvk5WGm4SAlrIFI08+98vA6L1WTyAq
W3+5QvCZbZGB3KFhh6jhwRZZaXgHMifWpaFiIrWyHsXtizHca6zUxviDSQlZmNDEZgrIZythD5tt
F8sdfSfNXrypw0NQcq1odLX4WKQ+EaICinotiRqjhsy4OTvffwwLKoIXipanNFIYBoMxMgRthvl9
/kJXaVtGNnxiJHTWl8jwT7GT6dqU2rLj7v/raLte16oqmQW4BI3QSzDeee/lWURpzFXHNivtx3xP
p4fQbl3vbp6xqqRLXvMK62zV+MbbBB7zdyLZbr8Xipmu2bmo6frDyF1G/auYd3iFZ7mSsR1M6lUZ
d48HddSad6s8JTwr8/Z+GseC/poLrmvijq8ayBh934J6lsOgcTexZKLj9ly4K2uwUlc4QeKtM2Lb
dXcScdcCBIlrpY5c10G2wFR9F/jwD+9ey1m9IZf0/rP+P93A8rFpzDrh6VxuR2lZ1Py/49XeaZzi
B8+KykMcwlzZtg9FhAD5DDl2Wk5OT2MHSa5CtuKMhnpQzR2WGPWHlQRsGomHOr9b1T9GWsu2sSSX
Z8IPZi8yvjvw+gqU+HcnDpuixixyY/HMJV8xDzYrKFfEoA6tcixf+X7nYyQilymUyWlpxUc80Vp9
xh7LdGX5OmDmpiV/xX4tRs3p7EQCc7QNu7p91/AUo8+7CYNUXzHEfbcQiidUTvL+aIpW2rxiZD+J
XftettFhmeawjQqQey15X/EctkmjkI/WsFFkz1Cd21ps34bGQrf3DXqs4Vsyyuchuv9RI++VkM69
E6eBokjcE5sq/Llj9V43zECrlC6tHXTe8fCnvvznc9qWmOElUFBkrngp0giCbcpy4XUCQtn5Ci8k
mGYStZG9Ounk5sK8r43WuZA+4KI0KZdki6su7ZvlKc9mgqfhovIGVLzuRegqYz9RehyI2dV8+9mK
ATSa3MUWhYiZRSCTw+6Gvj0usXayA60W7xk9kq8kMm6wglDNjEJF9fhM61wmN49WQG+dHvKbtP1U
y1Md1ldq9mA1GYb7dwC4hWQrceDGYXpjw2j4dqKgK56hPbqX1HD6lt8eWQDur35qwfGaV878a5kl
8C3KFlbI1FoK82rQG49xaIFIwzGF+qEFtzp9ucSj6vBh9fleEn/eFOBCRSSZWxpKV5c1aZq1tNJN
A66uJAgWK90C5DTMrxqlWrk7BDR3rebyreMKXkHOxTEIbB4b2IswN3qCDuBYCYoEwK8li7ZGE2pZ
q6+3RdacDWsP4rtrYs0r+oCGsX88Ti9T9F/D5ySIqmcnWNxlZwNXxOkm8dkGxIEw17lTCxhB0loh
GDxgTLHuztEHOHtGQY06Az23ZaYhtEkJrYWgb8llEwItYm5amMdHDzDoxXfQk8lnCxF37ihvWYpi
9MsEMFS5AEAnZJivjpS+zcZpGk6lmCTU+qRo5Aae53jKFLtLzq1G4vl9w623N8+KEuLiGaU0RQ9R
tck6Ncw+jRKUzeOkzr4squmfgLf5qR6egc0xdS/VltGVM+mZXCv+MTJkjDF7R42TLN0F7qCWsCp1
Jk4Xd6OgmWysTPIz0RWJwSrgv4gSAZ5mKNodCp3T+BxoR/hDrLbGowuNacVtzh1I58Q3wRvEbk/1
qJEyjqewzB5B1eT42iM2F3xoFvm/DiPXlIj85r/CW3oRas3pRPpWSvb6W/c2cCD4BuQYp3nLSUwh
l1u7zowZUBXXgX8yZDM4rYi+0iPl5bAPrfN5EFRhv9KMTPUZfI6NVzDpSTi3sFdUfUqvZtlkp5sg
b44KM87kxiICH2PMzZT2NTechHXaGbDNr/fa7Gglo3Rfgxol1EeK456KyLoV4V0EAXbVpk13mClh
7zQsVWa4Z9yP3xTA4R/4p4jZkGRGevzYtU9lU1iAQBvkZ4A0d+hJJdvRdlyBxNq0leXWRsomiSar
mqFsRQfldDGATONNI1OUx9qYfq3ydLAnZChAeJcuJx9OWrt8N9cMBHnfamKN9Tf2391b1oFTXstb
HBbzW2bXducOXKTdWl87f9Mm1xQoJXF2RJke37d10F8eRoIXzXLAvw8Bfz432v477JKUvJ/lcXaq
noJ8c/PER1qhVe62fhhaReZ11vag2jZ++vN6TkQyQRxN+JD8Ss2lCH5ABbMY6PuxWerWcanYF1X6
s+ojDh/5nD18K88n0gcm2oRJGv+NsbsHmBFTAkBecBBu1WqvgvtQQz8HcBkKm+uYvZ/2ECyQoVfz
t6OM5Vl2BLNi0GQEYI5b7k7YOYueNw7hMWEk0hUhBOMcqSfp96WikF9h6b5RP0ctFCqnSWQjAGWG
vDxuT10Z4QSHYQKxFgrOKTaBEfKndvKbx9gwKufG9H3tjsYp/zlTLwAbJkCgLCKV2eRLEGQsTeig
uIFOtx3SeRq390EkkvlAm09Mo56ezKoWri2reAs+Oe3BmrrGp801o6QpgxfwOnR3nh/27pWoGQex
wzb0x7b1Hyz4GKleWtetXlcwzPEIDhF+U3lJX14/Wjn2gXtyNFlqqSJAXqrM0xm29cVHz4UUoLdT
ru+MGjwDKyZShidTcUS7TgU4p9U/KtAxzrte8f7l6PO2ujbjiTU6ioeh9cr2iRxaai7PFghcSFNE
JJIQF5+C+ALO28PT/LxE+wa+8COgsoWKvOquQBPPLvRhfwjjcjpD72M5t8slSNCLY4PxFCYIVkf/
PP31Fk/6m7DXOjqvziv/oKi1GsTfD8jmsgrMAS34BWgTIAoEGJJE2KsT3jSY+WTcRrSNn8OYWsmE
LRlimWgjGHUyh/bqtMkeVovrc5nEJTaeSMJOTa/xQjg6Sx/on/+ZZ8hw6/3WwUKI46SetBNHpR2J
blbU9mT4lTQVxtViaaeibKqTBcc4ktMbHl+947llVYGcwwTYXnWSzhopG5LdSwSUpWdfTr6oVWLc
4kfSUxRXulYli+s4nT08HYmidXuhR+xQdX5F225py4LW6vAxD5oFAd7bl8CEd16mAuOqmwvcLyLF
tqMdvoqcce0wT1w88vBrddqOfV70BcagKT/dVWnInxb52q+c0an+cOJGCnyuS5PC9zevVc9jJybI
YXM2nnc2JXTarkmQX6oNRdAWZQSyClVGR655D0pvVsp8ELQEzMA1Fdj0Q1ckwK8drZFIuxX8h1Py
KYJmkGob0MNngkb5Ua71cBDLbAO67p7iGhQBa5XA1zvCDnfEv8+L/ialp8i2VGnTy9kGeDeDqBQ8
INnQtUbGAURzupV0uogvEYPPm8QLHynQQtWTpeTTZRCesXYZeAqITEzZwQCuvprdLBxT10KIPUz+
VxGulbRMoNfyvAu9H7tSvoFKnSDqVMrQy2tY8ah6R0za7sejKSjk3dwUHvfnVHWcQ70PnaUT5rZI
kYvW83/0+i6jCXPQgslQdAr3oYuvucWPzZeSC8591OZYXP6YOkc8KPxg21Epscf4l+xqJf30Dr38
Wy8sX5ZJC1HXN4LNYZJwUU2VZh288br8YUuSPsgjZuNt9s0wDVVxcFHZKmonlc4TssYJBYZefUct
0FndlFpM33jAPDSw1HpXraM5JfcDgob2VPXYxC3tGKRWAz/tZqoz756SKWaoUhDjvD+NdQDi7WcK
2ZCydiSWQU0DecuJoCchFelONMSwLcgjc6yf3rSxT4tA+D7lfONg/ZmO7NhgQeBWXVaUWaWMzFSe
Tvq+Jhqguxpi9SIG3XawYdFTr/u4r/0+i4yN2FfANw/YF+KCX9Sn7Uo3871oc57lIH0L4j3v+p5B
I3q2bdhvAAC32hB7oWYGNk5qlLy7qWf0X+iIvJBoAvvy9kRzZwsh6yLZRkOg5Coa47jz/L+vfhkR
b+kBNYZSIJTY+NMXNdd+w77TmSPQXrCa/1LAw++ssfTkyj71yidrjLnQlnOU4c1jZk2xdS+IVryr
s+RM2kdxmoKSfI3XQV92C0F6TDcIXT3qZ7ti5pGiMa4th2qMjxNM0Cp91IyDWs8B44Jtrv9KWMki
G8yavOlFJeQunrb00JiPjiAJqhxCBTkJouY5fZ1yFSFHRg0IT83oNMZ0SbW6EsFoPZBpbcLucO+I
BpZkVR16OIuiSteWUlKrYcgUq0EPdGmQjAi3fq+T3c4phYzh3s1uMj1NQV15i5OMUBG2LqzY6am/
yr9YLiJJoNZTcN6dVk8Mx4xiakqz+YaI4LULJk4VJiUWFGxMwwtcWZELgKcg+QFmmtP/lyKOtiSh
VnNavsvYxh9r1bFITkYSVo4cJDlp2LHTA2S1bKz5uep3n7mfGNPG03bYBNIcvq6E8lC9ezfsFgh2
FZY4nmwvnTTxQeit8gUVLXrpUADaLyIticlJBikDPOCRcV58y0717BxlbroQu35iYr29B6tPf9L7
1lD9pRraADTYmPFdqd92AnoNmQAYyheMOlfsWeeMceCJdkk0mWYEAB3qIOxbtjORvq1cr+Z94yOR
678euuPgiJXIKew9smiy6B7/13Lr1NIK637r7WWkzP1ARA4mMAvSFRIKY0z+dOmqYhLWha0jzN0x
/yV6Q7HCRt6jF0TnmANLILbBoiH6n4WZ9V11t5m8xFBJS26z3nmQao+K0cSacqQUx+XbifznOQsy
u2PxV6yK4CcSJXCnz5QKnMG3GaWK0U4rNHy0VEhsC7U1GbaWSVAfhBFG7eZLY4KyKOhIKiRlJdDD
F9vaSaVMvjJLvtordLOkSQc0QwhoxylM6Ln0Xzhuap5gdjz6iAh09mhKefse2ZbHYRj35IizKxnH
ofmcrEZ1F/BOz21jKtJhImiedVsxa0Mf+XDs77d75M4DHcz4X+8fNoPmwrzjrMz78oWKkK2nbpSv
S7N4X/GLX2i5mmsxxsrtkrFttGAzudyLVEAE09NsV0Y8N7jFc1Rr7SDoNyMaV5ITc7GsQJf4Ew6V
+JT9XZf5G8hBnh5LyGTd7A8heJF9VPtQxjIHAbZBNwNd6kBqpsklOZ3g0bDfCQoA2IUZuMz7hK0a
d7ZL27Pl5XD5oKHr0OQeVS4SBV3N6M8L7STb4Khlhiju59h/o+uF4Q8V8Mju5fRGnSv7tm3zFIfK
HXqN0HUFdXZVmK9jhTOzQGVAECSK/dv5qlJlehXzrYI7SEGal8NABCb5kJ1a7mQsVRggYgvBTfZs
iowng0yHns6RweY1wWEE/V2xHyuCJjF4xEj6MmWqiJRLXWbaPVjNPHjnnX0/Xo9xB5uMvo0d44Y3
+WvlznpTYl+/TKya2VBghbwr60idlFjaXkjmENAZLKsi2enS0QMCLxrBqZq1WNbyGputrFEtMFan
03pATlqxsxRLDko7Rlgu0zKJnFlRr6Q0IiZqfAX2IJVGrueqCgF3Gnny1z2+I6jGwBn1pTZ/MCOL
mv2SGi0HL4PC/NKloGHTHV/CvzMAt96OEqFHUs5X8xT6wrUoQV7HRvAOFBE+si7TKUnJLhOPIt39
1sQ9gHMQKrkYgWuPaaQPerJg22ccpWbv3atqugE7rPrZGvV+uAfzG8FSEhf6otKqD+o6FUGVghil
XrpYqF1jDItzZGDWNNywumLYqwO1f4BKIX0x24DLN3Do6YtPktaWXrZV3GL4xuVIwKMFbk1Vtdne
lz5PmZcHUyG349PVVF6b+koeLJnxpBwjQTJB0//jGrJBKXMPHpXkvN4poPlAP/CHkgo5vicNCGaH
QotNN2Qx9RbwIURPMO9vjgZTzXEV9KrJcUBsb41BETszUeTFd14i3JOXs0LdC3SPripd27v62EEM
1cQ75MARgn+woASsEevBNERYVhLUH62XKYyCB0b3mQ8mSL2ziPEw5GKHshHzpcO+M0pCHdfmmWWE
5yhKGOO/8ln6+54fl1lwTl88txIS26yuWIv5+DZjP0TTiAocw9h8qDl1mh+72nnMTF6tdR6TL8N9
sGvB4adPLPOQL79QG+Dq5n0xBiQNgvL4a0wK4PNRcRRtNO4xrtS3WBNwPZFBGWtsD80FX/2PLTGd
J0/5/ASbM7lWOihDZT4oOr1Q/JImzv2grBjhqVPapuFdk/FkZ7ZcoIgV48kaxzbLq0CdfvF77xDh
lgHe4Api6mgi1UoTrAZ7cntgCSEe9YA/9Wj+YkmhTHWk9k1Lsstzfp7EWiia6gVdf4gutXw8WOBp
lKeeHAxPDqJPBkIcMhZnOhQZg1QLyTH7NgFI8NAPZLcYLg15E6N9H0FekfYGE60de2KMuXlo75Nw
GhNI21X9sFzfYloXDmZL7kS6iPxba4iv4ysX3yiKHEFyGGVNCKaeacanAbg+fE0Eyfop8dgUeaV6
vR4AE1whkGL/RQNtGmxG+yMdCeX7jAJHmDpZvvu+TMDgBaq3BweMhVZtpuDjTNLJmqHIse1dJT9E
7hD26sD57gGSk41qr94EO8zLgIRoGKftJzM3H33G7+lLE6XrMrZpS+KHs8rjIxjYtbQJhWWtWDRr
oPTzX9ltZzE5O9dRh6Xvwhpm5ibbpLGfFXN33+/Epq3vn8PZSBn4mcx2A7Xo4spyH08AluSX4twf
F7ETaSmYFb2EuBAFof/f1AddgjgTdUUonsoFj8lLfgOHMcUI3apNdchkkshUypdWpBXASn5hpuH8
qhNFqB/eqCI07UKxNl+X+VGlO4KTEDsO94VD0nYlEuYoMnXT11dVRKmZnd8ausSnZtDp2k73Qem7
LLcQi5bBigPx/PgehPc8Bny+vO7a+GhCE1Ujwy/A5U3opR4mRjzz9Crgp8ZgDDS6LPUj6yGBC/Vm
o4gPjZq3lInZ7j99Fx7nBeRysMnYhmwR2xvOfgnwbswkIoLN+im/Pdcfka8Tobb3E/CenevVnHP1
kEjUXn12qYgMYx2QMF1aPEfKC76gEirIcAOXLzwqS48LaASjgbMFj0JWzcVXhUifZbIMxmnt5nJ4
hwVwSAKN1wcC0i4y2+Z7Re8puQSALA9Cnz80ja8TkfKDMI8gm5eJrOnQxO2KPfaBSwmYfdXJVXSL
6ce/AZ9tkkPWeysZDjapsYs40Qndvd5AAFY43NkX6vQ9FgAYSeadqr0UgY3uFhZHypZuQKbeG76h
Dsf1bk6QfZmxLGCoAM1PNug4AsuD2yR0z4dDGclZwDqPRkntZYr8HaLBnUa22AZXC0eCpPddXLqi
FsFmW00f7WcS2dM5PfPAVNVseC9+7PDhKKqBp3eEcmtd2XweUJWbqZwLgT5QIPM7KZ4S/kuv7piG
2fbms+Phf1o+jOINFIy5dbsTZQLqsMP1YZLBQSGWUGY5n8N42XpVSMvy5JfDerTwo7uS9XCaEp58
3+jI0emCXNOJhLrqZM2iuW52uOp+l7j44LrKiPABax12aLwdGL6rEdeTG4jnUOphynb0Mbe2nRaf
p4z65OKOfZD8h7xzC2dd6IM21H9wINA+TwLKhYB6yjt62HEnYdSIbFwaxpORBXeEeRcR68TKAUfB
WrR4R3VYUnm9cfC6gnOB4zKY4zbKp/KEdVcoh+C9gQLE628tZP8Nmzx9+x2rlyg8js1HMzQ72CfG
QyfstLNNweiKfHupTi/Ep/3srvKh0Jw0XO1zPVf/3e8ou18muLu0ihPcZMZH6j09zHWXuNslGOHz
vPYUuTgUuXv7++XTAMxemCrJqfV9rXhyi3DevV+kG3zSEWDchO5Tt0fg3gKCWryjIqsaXuxKv7M2
BKvrGF/PreFVI/XdInSO2K3TkfsrARPJ/gL2nQTyZ7xlEvBW/24tzVfJ7OSnkwqFvyXTvLzNbwuf
cXnHAITP0vo1OsmNmx+3RwtVYwlTQuRFmYShP3chk2OBrtiwNUXqsoKfXUk4ZklbkxE9E2OBS2nY
huHX8EYKWKD8u/0zxbgD1faskHq2Gols7tmIJdp7qzxB0SBD934kiGf4teC0V9HioR3f2D7bOjOT
Hks8CxXAuhZtHIUVWa2Ic86bGeCI0vgqLdSX0xRmoxApbltGfasF/NxQwoqZ/LRs+L515vfS9xFj
NnZH3gnEf7pj73ZQPGlJ85c7X3Mr83AELJiLSfhsWS1OgAjviKJRUwVtPdKz9N2cqKgaDAQ1S0VQ
SGzuwSZwRzUe3gDwRrjqDuXwji5uRY71kqNYYxDR0amTc2p6uIYlQTnl5Jge6V1s1kWErDvr70Y7
Iqixi4Pmy1uWBSqinDMNni1cV2MU4V9t99clsXaLZaGaw6CjBj3wWws4eEo4UGgU6n02JAc6xnE4
Ca4ct53ancdbMotmTj4HdgnL/uK00isGyYE/YwEzVG+rkcemtzGrer0oBy5aVSAFLZlqVVjYOCfO
M4wRm7CvN6fCGfHyNE+kav0CgqvGtSd9SUpWVb3UssSICg1NSQVv83VzYoZaFjV/cpax6nOK2S4S
6b/2XfQz4iKaulZ8lzQfv18iChNOdu0liVJcUHPUnUDHHrs//T352lWkOb1hfaZQLdlMX5kPWRql
oYkAn32gjJmR5T6LCvJLpOc3wDstNZsFOBSQmgBM6xXy5rb4IOqRBAB6ATccOEnqiiMS7MZrYq/1
wEguTu7lSMHuMxykSNNxxtqsaY1GWRFe0poyP7wOn02ZqxrMt0dOTdJ/wyCQdDe85J1GHuFqW0Mm
bBYRJF2K8JPiYzmjp8oneuk/d+3268Afit7gpWDr8Dd/ZYCyHyLL7GAFfeAh1+qPYlp4IALabozF
ijHEgPNVaaEHjmbkczLlTaHTUkAGG/FTmSot2lIXhDziAiZiPktLYqIdU5P+c+xR6Motze5BjByC
q9qFTqHrOnVl4GTfJLcdSkKd3wmYS8bnXPzBS95m3wNFbsWDbSHLv1tr52ClS5mQZK2upT5fUzDz
2AlAw8Rs8J2k4EH7Abx+ZMcooKfM6kikmaShj2AatOG0duRqL+U6n0+EOOg5KFiBJ1PsSQfd36xf
Yp+F8xC0x4hzBV1FJUVnO6CNJ2Q1alEUgTEleA2PRSNO4J7FOr/XN3QSmH7hxuoVE8t3HEer1k5v
r2XL/wGXU+XzsfWCwSELdddTJqK4P7UgXhHdWovgFNVl/GCVlR+sprczDS7XKEWndhlnLXQAJqxr
h0efWgJPQ3zlp0GVYGu+woIGBCAN5YMjuSgJEDpQIB+jL1Dx0Mf/EAMNig+Y++CLR6lLc70r5cUA
ic39gw+K08kDVqsK41d1B2gMnd1aDASvlvpPEe3wWoIDhr78gANOZIQuGlOd/UV0jiyGYB20KgDf
WlWC7wbdt+3KndTQXVGq1EykfFczCC0LzXj11z2GUpH/LlJmEoUWp5FmfhWt7KJ6MqfFPj0tHXUJ
pKgp12wgLaHTwB9sF8uyMrPvuxr0nJLEQdCXSdWxHttOM48/z2Vge9BYKobPQH5CfpnFaZydZ6b9
9rs6SalMnQnV+QVO2o3/dgqQ6PfoLmbWSDlDi3t55k5tu5CwwLJNjZqA3Aauv9cTnf3Z3/3RsfPs
CgFMFoJlMkwB+K1VGWcVp59jdET4OQaXPkOzHSzguL9prI4Jdgu1fsuS+uKeZVJ8+1ihjGDe4WWQ
tb9Bums4iLDlJTs6/EwtogCUFnqu4nuDxXNuI3iyL9ojc+8Jxe4yyabQ+kiJg8cdQACKdnM1UtQh
oQMVu1uDGVX0DAWRT0FCHvYl8pCUnTJdBVZsVD4KvW96J5twzz8H4gtB+jRyG6z251usccqPh0Oh
mvtuNYH7sBe9BrhdnoeCYmHppa8UTGLlh8cD9DTcPgAtl9Er3XgXSE7vqgwEG1GP2CqsXfGZtVsv
uraoPTq8SeDjXnLKQHM5K/+AqxzXX4p6JA1ZORATAFlCsbkAW8wWMxIHSICiBkdlnj5qo84W/3hL
qUU6p+mss0VlHi/IwNCjQ6AW+s5DF5qqMuIT3uiUgWWMt6cTmiVRqCHAiScbUqOeJFYWP/Lgl2kl
FHJLhQgFPXVo+4w34KgGYePQRfk3daAkJcObc55lb5qAMc/B9JXSbMyiZIOWYumCp+soIvT/HFcb
RRvMe+ji16uDUK6Es/aIHmGIIR0C+g/a9rbDUJswFXd5jSqCiK55FrJ9yUCrOw9Cs46Nmrh68GTg
HvCna+oWAKQpmIw/mJmmiHnV0pJRAEXYalHdp1bLzuMZ+vnDFAxk06IuM+wNkS8Gh5Brb+15JwCj
9cZiD1b8OH7V9YgrKC0zW+QFEs3EBspyPa3O/D3jf5DIvoSyuA0Z32fy7B5+YRIhMOchISy4Z8XO
KIeUZZlIHZ9g1kGs26QN5XVQtBqs33rNk0kfASe5m75kD28s0kmaDe1jSQsTkxkLMZ12USrqKoer
q/1TcNS0mUdxot5IxfrT+FJweLKRppvUJhs7GhbV9fiw521WCeeRhPlUx3joGwY2Ez92xW1wFdtN
aEvI8AnssoKx3g30KlfARyhfEFTXGoUy2QIJLvoRpEdFT9AO5LGyfLvMgZHf+o31iakJQN8V9k3p
hv5AP/rNDDKMoGa9L6rt9t46dxP7mLKGEVD2mQ979kg6wkytC6yOmUerpu5qPcMKNtSiaq/snnhx
siML82NQwR5wwT2aUhE484su3+DgmRIauYp+C1XvlRgxV/2iohJ5gJhBwlZtAjstqAzFnWqP9Z1M
TXg4eknFm1nOxeUptWbd+ldWwMau/XyEkpDnDtf99uilqL626tbTo0SAt1/jD9pwdu47Qfq2Ilaf
4aBJhd9MTj5Y27r09VRiWIureLIT+n5RogLJ7u7ZCtO1oz6jK6eDVDRW/x5+avbjEwm1aHSqgpFq
FnjqiwqMo3kBsuRrOfVXhjlfpd7FOyPqcgkBVSrpDSe0Xax4sKzZUreHWekAMxjIQNEP+NmoW1D3
991X0nsloWy11syLAnIpVKTqVT10k2aG0maBEKvEFF0LsleQThM6ZbvIkgknoLu4KAM0TT9zikat
9Ea0QHHFds007rZfwDmzsORjbMhfO0P8B9ae8MuwYUYafEddGxw9Xwpxr096Wdg7pZ283g2bLmJp
tOqQMU4bMsJjH76VGkYl6udHZKToscHuqp3mKugRSMiHAWg40QCII5Glz9adPBmlWhyU4k8TmTDa
9qxHEA0ExjyMf6qUpbVPsx09BVHfsZ2oKWAf5ih/g7GoZQlnWV89H+KEH9E4sUyvbdAeTWET5ctN
g+ZD4jlWOeEiqTeJk0lUGfFh3b505z/zspZx7OQnwTxuagRYhtzGn/6tIhKYPn6x7tZ/w1Qjq+8t
SxYby676BfUTczjSoUn0RUeTaD9D3Vx8tNQ0D67Mottl6xmGvMPyJ+nagiwaOfAbzKynH6ilFnrK
52VsvGEr+utP0FGNwPNfNNmvnbk5QYHFI+VnxGQt8vZS6JDwVoGEFd0YxtvNo9EcquOMqNTBFIo2
jMrOrTT163R71Z6Pdn2h4BmirnMoW7fqi1nqBWiZ5Lek9NZ/tY7KNMJvJmLpAfLvlXDsmFIDL4Ve
t15sP1MPFhg9WoM9TPtOskabeWRDU63mNtAGFXL5+ZE2GpMz5BjVPcfjbvLbLNvDjZWKpkmRC2+O
Nm9qBcDA7X6Un3NRzDDK/cxiRr2jpFZSXsX5lsAelQU6agAdpX9sm/BhK5w8AsyZwwUIxEB/hxvh
b3nMKe4PsjQw0hnXfqkqaKkEFu1fwdC14TiGmGL8/DTXTZnFHEQyYWaicOC3EGV8Y/HI/X88l6oy
UNiwhaKLApJsibP+c2IR30H+QRkD0E9jiIkRAcQ5o/YI7nQkT67gsCuxKNQNR6Kxkvov0h4gmuiI
p8DSFEfLFHOru2wbgy1fRWIubwufgpz/wXLV5poE1vcMmSMHgQA1qweO38rSb37ulTEAEuczz9fD
g4uKR9w0aDIapUk/stHI/aOR9ALGSrx7R/FUV1L17Uo6A9nRXo518o4F4hR4ySE1FTDKhcLw9E7R
ANOHPz8vqg0tqP82WPNCH2Tw7phyPb+P0izHcYeQ615fYZDRBQN41bqThZMEyDOp2JcT0gV6CLN8
UOhZoYcxsxOaOYaLVvVVBABWcOr7f1OzaVvoUukT4bu+Zm2+4jBldoguWctGuxNyEax21k1TyDrV
bPE8OPyM69dqHr5nKGXXaSD+hvThDowX3OMgxFWUNQ4KIZue1xY5d8RUZaVOz3oVBY0zQ30UjVDd
wRvbhoflDGEW8CNTxCj+il9HI5DAWBjZw/oR4Dn7o1JImz++zSrH25o0Sat/hFv2/eZUjWhxfnah
bfQPfxVbld+McaGAPpyDffLJyktQwBpIjVPI3S9BYh6ZmZC2trS+LClKSiuFaUia4GDgsIJ9T+rM
C6Fhrx05RBZfSC12L5GZ22hBSJhI61SkG4fp9mt5XwbX6xGsjSPb3e3fHmmuyyMoAMe0TlHaLWVv
brXwwSp5hoVTHAh3dQtGglPlwmWtf0mm4bpck/6rxWZoWScChOQsVzgG/sXYpYx9xZiJQb5Wyeby
epfPS+IQ5IXFi2+IydcAsnMBI6dNGNbfRLoF22iCLxvUEtqmPoouzahkNmoGYKVLHCuls2bGP13d
VH2oiXiCPju936MvYvWMTfujOtoDCtYGeILGHICnubwkW40mcbFTUF8iPjFSAwji2mJmKf8lBBte
1inqCMgUvIJHF/uZp4fTMGkZIfnHQvBGHbx7RXGN7ILNWQz8aNvX79habNgyjgQreBtvD1D+pAID
eNqWm3eNUruy8GWDuppUQJqya8nRB5FAG7Z/gfLWEK0Mrk8jFyJxxmoxyZUp6WNLIWGvkqptknyH
XbrrVXi436f9XCXFer3WJoTo2lp1clvWTzIpPh84K9TRYDclKXv0oRipOkkS/XDrnPtmTom4hMj7
T/zXR2aKlxELrHxNLA/e994ciIWkA3OuQomwp+fH7iWfkqno2tCUA7maBhvokksg5sUmIlxle82G
hJNeb9ihPAFqNwPhom86i3MRjBZYOG7Q2eUMdVoyqJUBYHq7hMMMtoUFPWmyAxQXJfuF2pGAxSwp
nYoIpcUAyrZgJGVmLywN+LLYQcVktk7FRJTqtLtz5IEiN5Nkw1b/tORGlF8Vl6ORhMGvUiwPpovV
H3pP/5joztGZtyXeDUDa4FWYlboIfXY0iLuYQTz1daduZPeKdoqZF+pGPLLiYIzCp0yGyc/3D1aE
ye/Xn2CU8149pnc7BTezXS3w+jGsVV2jJLNyvf3fGx3Z4WgFbsFROu6P1q64wn1gNB2VC8zEcYAB
ooESwC9B4X64jqeZ0SvFPQt0ZDd8YPpHuz4v2Tf86q1avoCWfglhOCBib8v0/XGQtcaiZaEEyJDP
+gGWpNulrRwQa1xT3tPL6BBCwbi48Uipx1zQ0S5ClDqqYHk2lbqcjeTsC9p7KryGhPTgFUrxePVb
zohspK2EBSjM2aLjS9QBMlL6bJ38es/aZA/qSWOVY9TOzdFHgNMMgs2wFkTULdGMborO3Tjpdqv7
PTbYh9AavZLPEr7+AftUaBRab1VY/Q1bCsDLBsATJliGDnLgmBLmiZW6dy0YpEOjb8vDCcgkr3u4
a04HCLD82YKEU9kpfc673SUJzxtrK1dHXo9KwcWR8nsdHQyhV7EpprSka7DBzzvAwasu1lekR88b
kzvVvqnr5ia8wZnnWbxZTzeKd7l1SrGu/c7ZPbWQ+BUMau30HlcLMt8tFp8hSiQSk6m/Vqfzwoi/
ZKu6ew+B4EMZeiZw0c6CO9otqi3W9Rtht0aUvC83wzifl8BNLko2+wfL1KFi66uJg0zpUprxPAP3
VYyjkCUcF3drVp6h/Fe6rwv96RtGY4sS0u+ndEIj8OwgxpqKogKl5SxXO5iE3gwsUtUdS/inkGeT
q2jbFzjkL0H6TyWzngNezwG+f1NuXUZoV/JPkUsCoGMoqYibA//byn/70WBVHHqJeABh6YtniLr4
iitd5LSxaLkch0mq07Ysj3vaZ6Mhgibl8nKukLZa+f8MFiwLNNkxCpzaG6N4qOXFUTl8paLkpWHw
N/CcNE5edzfPxs6c7xf2J7irZ3xz6eNxp7/OVY8ymFq3Np6O5TFjiK8BY8+9nutEuiLfFK2BI7/v
4BUwlMzZnWlZIlgjhf38onKdaBXYrk7pbfmgB7Hj/XFyuXfOsm6dvqVwM9bJoDkjaJ/WRmpSGYdv
xkqWr+a+XsTD12oc8sSmRsxzV1D5f+sI/NFhs6Gv3KAPqgdpKAew2RUNlypHjdKPr0Wi60Mywhp/
xMIXDuEY5e1a5ImbMDh/eBKQwkdnwHeHcKQISA0NWvGgpjoeWZc5yWBkvVfTdjgUD80mDcjkpweJ
M7SaNn5nMbjFxT0tLqbheA4biQog9YkNbuvyMeW6nxyRCBveTbaOglohVB7XoepPQwWeTuVUMk9L
jXc3KMYeYuzo6gGC1MRnwjtR2Hyp5WFDTMsjZ05uIZfCVoZow5154F50q+bWpWckJuz4I71XvKlL
BD12xxZDtw6hqZ0yzVuB239d1c8v+z+hNNVShdNF47K6ku2caEMKZwvnTcHyq5mzods68IErlNSh
7BryAX503KMPDT2peCD2gqSU0i3q2p0fSEkSrhUNLgoBU/PWO/RQHrhkDDg3I6iY5mbER1hETQV8
np7LH/Xoi1K9nV+TABcNQSIDlYrCpyCIJuEuRda0QoPnuxxBCmDGo1ZNANxU4qd+f6kCKWTRmiF+
uza7REnB3dA5SHlybhh8Cg+yWUjon2arwFPipYcQAPZr+fldhlxilJa6Ahg09XJGMIUKev0frba9
Aj9J1R+EfX1c9LUgAQwDLtLQTdnWHAMyGWWWKOipOlMW5CCyUHHGO7bykCEv+m2HXgoIo3QKaibU
7/CUDBq6YSss8XArw5AFT2pyp/OeSC41isDrCPrF43X1JP9gvyQgsgNqW8CF8tqd+KeOHGS2r0J8
QbTvHxy8CAeK1Rbb5CExB5oVwTgN3pYbz5iwA7RatiurCyiePk4IkR80/+KCGt1e9aTSmbp0x3F+
Jkc8qPRfsdUvyC3GIe1j+A5rTdJ/9dTDQ3aNiRGEHSPPzI3CsIt2XWiBFfF+0ezt1OiyNtFoY2qd
wCTT2pGQz5nIV/hNsHp+ZckIUCNIcMyoMw3TgOdUy2vae5N4DX0tf/1l1qM2quQUbTDblYKY/8FU
TiYt+qYyrf1NCmaBIG+FgZgGYm4xb5Vs9C9GonzCgQp6I1zdGdh94jIqaLNKUgpMPr5uvXy9aqwH
FsaGT0OBU3siiTFfa9SvL3PVYUF27PuULUNxUuwPaDF8czoQC9DCPnS25kCuLKjN1ZXqmz8yI5yx
6aLILlstWA1x116zw7fTgmCbCXl+naMBLyUB7yU2bMurEMX2dZuWJuiqUHVNZOFVbqHsehbgzl9i
+fDFbt1DlG/iHdPJT9D2hMlZBGXK7v9D9jMpOlkiIk9+s2Y3I114uMYcVXnuqnZtM6NUBLhM1TFm
LKt/12aBl4LxVZoxEgxPz5vgdVIJvq1myQBeuMipuoVHp+iRaNcUnbzu/eQt4sFSLcWsG/zATMU7
hvt4q/RCa8IRrCSR7gJOUB4M0Ix15QVmiX2FUAnpm8aWah0/ymOSDxNxi6na/Wszow/HPq6B7kLa
JWt1bRuaC8eiIQsgzhWx2y3hlgPBkkXM/ziTOg+9z8/FkiY6HBT++iKlCkgpAitX6/uOvKsCj72s
g+EuXM/uJmB2oafyEp01GHefZm1i8lV6mTJgB+vTAd3ybnLM3U1GNmoOVgJCQufiVW1gVeYt+OHE
LhFEnsOGFRUUY0tcvyubGMEhD4F2/+bcE56iv/uOWC2udbtKpIbLixr3s+r6K7Y4OK95GS/aHf6t
JS5tJeL31aVZ42rSbnJiHkOLk4VvgtjGSGkFpDkSm182rPwb//n4RyR/+CoANtazmsMp2mnHZ/oe
q/A0/Ls9EcL7jyFw+m2RW2MzdROXi1MgjSHXERUDeAUJSNGLtNp2Ai5fKpIeGGiamKGg4OuUfDYw
XdTXrZBU5LX/9SM8/icjH642AJkwUZzF+D9I2u531YQoUuEYFOLgR3pxmJEjTgZdarOuLJj4/NTh
lFfEmp+ZSlxGEHf97tSPmk2qp9E3+/RTLQGWCwQsR+dBuldtwQBF1nSFHGeAORVpsheiRrrpbWfF
uO9qah5RT7lD1y6rmUX/e4fqB46mm2FFeYcyAHayRyflSSqWDqGxVlQU0ExhEHZOmumuB0yK0NC1
n9FpgGeoW8L9LXqbSTPZXTekkf7ICadDYIRv/rtuXlDlc/lq+SA/ZHdCdTGuLOvnaLwONZW8KlrV
TEsnyfD06wzU06cEmkw+LM3XuCEsywejCAo5/R+aKFJclnjAvSdhKjM9WAvBRFnKkHkJvEhC9FDU
Gcq21WonKF4Y8pvVuf6+JsTiz5SeirzCliKIqNuISjVjtOMm2ZYN8OS1c992u1cOsmTKlUAQuGLA
ZSa22R+C4wD2YhnttzL+gQ575BPPI4U8UYq45DertA1sHwJ6btD+PQC4k/pHWbIhCUUhPXN81PTS
TbMrv/bH250rxLhRan9hevCjKAQKaEPERBak1yj9xonV/wEcl9NSKYCNFsYKefanu194H2xpa017
2+RbsnA0tfU66FQ7grcp+/qqn3oaNKRAW4mbgoOTT3jAR9ACTn3e46HaODmy3CwJdMP0JEPQEAdV
M3xsN/Wvdj1i927fT3p7JfSs7by+NnbvSqqJPr7whOUoB2NhPn2cmWmTpGgfi+UcnmAnxqOmjf3X
myABaRvBJJT5FpZ7Dv94oEQd9xQc99ZRsPsO0Zbvj0iYLmwmpQfWg5aMKtAmNmzY5SbcI18bLrla
nixRy73KI7Uk5xlhV2K9u5ei1uwQr0HO2Cf4CLpBUUY2wcFsj8U6HAeTi+QHhEBFTZOHEtaleF4X
8dGBOK7fIa/F97eFLFyp0oviHxLy8CPglMmJlLMNM6idA1njDsoGvjrb85Q34z5Ng/EoIeeKiM4f
y50peEY1ctgWADyEEyAR4NUVG+ORk8yXSq/K/zSDYAp55CROLCJx3bVc/yTFxXXUPsmo3Ai/Ezhr
DQ12KNulft4dWX4dHxQBJayUx4wBBuvR8Cj60xt7NMFwUXhKcBOSdZvkjGa/wmmmjYKbmtBkdCng
RDgaQSXD+LINnw70JRbhQSfsJbJ/+h1Xg2LvOvx/4BwfZEVQzkq/UD8ajdWnFIk05YHDg5HQ9jwW
0f2S+WvlSJ1eXGmYSh2U8wx4WAlmStJ/moaVeuIFxVcEaRvc1NUhE6fh0gs+ExbaYRKBsqS1Xt7F
hpjoOKqgOd6tONWAxKUjfMi0h9jV2RjCstkQAiNsH3pmtNohCOwea8ube7yVE1r/0S5UlH85nNb1
WxCdvc+N3XJQtGHX3Aj739aNKoFwK6hvLlRSZq+QD2aibqumoFXPI4VF4Ecp9aeEkFZX1tz5lrCx
rH9kXhKAelBOthc64/s9N0rvyvEmgFJ7fZn3l+T5K5TREWQ8wbjNZsbcI1YHohnlnEnzZxDtavvv
gzZrIKks1lXvck8j/QK9jfCEuDTDuGn77pGish4cROmT5TiV8JbQUIRQwQIDD5CFALxKgTiZ7c6R
kAR33f3VKt2rEnqZVspaV7U4i0oJAPQjk41MsiAj/LUfKzIlYKjL7oFftaPihr+GR6I23R4pbIiF
LO6t7qC5Z8N+2BmQIwrCTHjripEsgO/Pv7lz17elTq7Lf6qWnTmu2sUp8Oj5u4a1t1cdNiZ6+G/7
GtL5SBOwgS29dd/ex0+kp/smgwh6qqgfy+xFjEL8Zdt48rbg0yzkswFXX7aND48IC/R7sXaAEXXH
6SxryMRCKIW36ZSsjlh68vEkxSh4X+hEwwOtK1G61Rn94IWkEo50IG+5uYXz+wGAxB0VOvtffGlL
PHBGf6nN2GtbwR/9sxDnwTYuJhu2JWjp5r78cFjPann0Bc0UsZswgpSp80uH1lvMxvvSPjaBwEPN
0JKslKDhybfH/PP8H/1fMW2WwpC/dObnkOZreEeBlnvjoWivB4KAjc64/nNB8g+hylBqA6jbMkzl
Ml7pvDCtN6lHT99iAsgghZLo7nKucbzVqSExujWr6J5VKJH51g7a3Faq4BqEkLY3AHw8MDOcHwrR
CQv03RDCWNAtG1ZrqektaGCvpSAY1aH0aX2qoJHqSWWmhqS2l4uf59Tqs6NvgxM9w5nR3puy3n6S
j6pOoTmDGGyRWti+h2iu8dNYwbWA6a+Cbvzkx1Hw3F8Lqhm6uqSk98EvMIl/LBMOiqZ+/1BCmrJm
WlllJ4rTBRJMna8Z2JRmVlDjGFco7DZlBCITbddh3gLeHjoUJbtrQrl76cWSuY6YfQfPqJZm6/Pp
gpjP2tETIPaRjNezTHegtUyRZsFkxiDeepvLg0ACjdOGNdMqHmGup6XvNibkvo0vYdoGOx4W97Y0
sS9EVBZHAepLqoUIDR5ukxafdFvmse24XOL83GYEzfrdCjDII7HN2od80j2okrXp37XEBjAReybr
btpSO+oXyVsetTUZoyvKM9ctsoa1jmk0mqvBtl5X4tA2xY5CpVn/BG7CjboATU+XEMnOBX1BivLa
eigErfQs0YMwMB/4/oVOm9T/biqbKVJ4rT+uUqzIPecGYADFdz/ZOitw7WaA73ta4nEVXSmZGod3
t11um5yjgZCO6uQws46Xc3r8TheF5gkdnelcpoaFlPx0ErgPEp/AFodRoEUy1u176+Ch4fCgcUQv
tTGq+cnp3DdE7m5bBWXqRZkcCPuRxjeHOOElBcVF0dX5nwZxoVdNrjvxbjMXCWuqhMRAdSTkaAPd
tNh8k9bB9AG804dq8g1TxU+M+ytVlgK2YicS98z4i8qXYGjEajvaVGLzEUQfPOgZhPc3RXXcp8MB
mptJtAw3ZTQqP3X/rb2RQPN1oT7LQf7hGQ0VHdibts/e/kD72+9SF2NKRrvmg5+PSXzgCltUV6H8
LryeGVeDULvA//gs+L++4xwcKUIfiyB+6W5OXQU+7Zkeo72OnH+TTYV2gF36lq3iveqqA/uZhHfe
BRQ7bPxIf5zs3UyWlvAJhFB/a2OUy1q0SX8quXBKLGCQ/N0cI6PBujhg4LC2MppZ0pK38Qcn3quz
6ngayRr+TqgxLXGTG0hD0G/Kq/I2E/9udGr1XorXn1f/6k6+JqCKrNzIzK5svvFkp5uxQ0HzDsn5
cUZIyoJYTm3pmrUvBbGLaILqG3YNGN56U3a510joxsv3KZ5sO3AVHxu23q6BLeKtB1Gh/is8ipgD
zDIIvSgtYmq96Galx2z91K6Z5iq5cmzXijykrJI1D7KrK3XXICxlSujpHGitxxPuNUoQpsToDCpq
/y/eMct1MuuDfjFwT4cU0bs/tvMQdebQ1XN/F9TSKpOKaPdbo4GC4zAKRoqqKR62uIs4YFw8qj9p
ViP6JCWcx4Q2qopIteY+4NuaGEeqpdzt0dBCoE++c8oPiISA0/Dua6Ep0KwtsSHRWlwUGz7hSVau
v0nSCnr3OuqUHp+u/clnnc+iuK3DLUpHtsTOO/cf+mWAphcF/FOk9KFmKZ4HZOgO9EppmN6N1GVQ
92r86DcyyVvwdKnpYWh1NQO2gpxNy2yoBIExsvN2PhDdLgh7uPdRSrkhk2IOprQK3cn3gcN2seGA
dOAT8Bp0bEOI6obLomOAFW5xJH+ckeMp1pUisJfHeb9Z39kbLwv1fLq+0EBpgR89oWWZ+56a3Yoz
rEm5CGdBNPvQyKBB5yZ9rpM76LEXae7OYLy72UVxE3/rRKy6J/+X3xUlvgwarLnmVjYXBPESoMez
JCZWQbzwJ8FX5frSnW4ENS5fRtGzJBnMoNC0Ktx2YECbqJYgiv1FTJ6CyigeUol5miYwSrCwUmfX
TImzvsX8w/3+YB3VMpBq3iaB4o8x/6NtZl+4PW4+i+ckdW0vLZmsjC4LTOl2kXcBarfuhIQGXaoe
1m/SVDPj2zeI39dCwB6YyXH4cwibpus0iKykWK41Zl/xOteFmUzhSpMGBLExMqyA5y+luCiID2vA
I9vOIiluM0H1+4cDYOxP+K9eeifdXFrqHSExWs5M1Uv3vRBveL3dxIjpilmuqz8D+S15wkLWNyRV
1Xb3CGhvRdlXLgQV5P1NO9LTKtzkETl/10YhtTlLNiQF/QPHuMWRaVUPx00BOCf3667us7fWIWrQ
7LcOlhaHlhw7wl8SAjEjfI3o8XUR3mC36+AAocdCMUnfgQ758JBMsuZBbUeNk4nleYX4QQi8r4bg
m4lPczChpZU1UDe+gHzY7cjMMcU+wvS+HddyJtPiaFV+4jGbbne44gcFJ0Zm3rI7lN98vUD/x9Uo
aCmrlrcKEbl0jEVnd1Z8jP4kZMSE8kEbgx+YYklD1m9qHtWJV1UGHkBmXa8kCCsQ3iTeeMPaVnQX
I6vhxS8SB4qFy/JmhB8RaRFdoH5/CYYyQOnmvRvkjzBZA8EmdgsUmcXJm9vChX/LfFiHz0proXRo
qPlrF9H3fAxX0V/QfvjfhERrcUxUNcox68B6b/JO0fMLCF8lAbcOZhtEC6AA+M6wsOjA4nUX6nPK
4WAooZa/1h4glG2chmYtDL0tGhy0qs3C3RyzHzt2P5yeP8SEdBFhtskxnS0dE0CYSqP9cCXufCaL
GAIYP5Sb2LQ2w1w+7iO+FyWWYUjaQQ1xtHtA4Rt5iZDTNkj+ZikbPoD7mhwiW3uaxGZPDxFbFsXu
9XNNXos75VjkckR9tG5XXvl2QfubjkBWaoDVIon4rGFdEXj79lrb8Em0MTHsSWvZz9MiRX8glXKw
pBmPIBSxDLC+v+8EeHyVblnnn+mg9b2S07qp/YZ2LcQI3SF63WBrmsxj/Exqn5bTfN1cXMqluAMU
WBGFkjewvSn/sSch7mGm3PGccva0sW0yyVB9jo3n4Cn25hbrHVKNeLhxBXzMEfv8cmBLSA2+f7Rg
9lksZdx1CJXCgKaHLkXwlQRW3hjPqEZSlV7Ws1Z/r9/r9vhK2I/l5JluerFq2eO0Q79bU3Krzmqt
Ubr4E0UHfJXUcmuJGGzpSUtLsOUgdnBRvvpk1Ag4gEfYL01JNB0ohrAPN1I8kVTMfSBm2OASA1S5
fmiaeKu5U6HEiAAw0Wn8e0oektNMSus4x4CYdx7ATfQwg1RsElsREDCsHb10DuW+axBUv7mlVuK3
+Zjb+lfQt2m0sLR189IZ/peg+MdYaAq86cao9LnraYneyD7eVj3ZM5wRLohRMdghwc/LHxLiZksv
czmYBTYAyd49YUEvP+WINsKhjL+2kxLdEt2tNVbJb3fmIrBQcn4Jbyh5QlBMjmQvPBaUmT6oT3nT
HzOsviuI93i2o0oi6wjnvmAPZv/8fQxM7ra3nh22yX334f1Skj3HT5CUrN1wFlNeA4+cLqmWMScs
0l3XTA3n6d94FBb8Xg1Q57K4hYpIDmNf294/WxcmxzkoV3pOHOBmA76P4kwUC6/NXQw+xd2p6S2d
5W7UCbb+Z1DktCRzU/dUY1QHg6ppxCTpq7DjcnOva7tyA4CpUJpIfkXWdw/hvmLqNdGDL8CmQzvM
GRNDlLjAIFaXNpvPrIMW1NI4q4ZdkfRX65zk3moXLKWnVN2MCOBH6lcWGn6mi+P2gZ8QtDFAkPXq
+mGIPXzApQ/v54JRocMRxVsK2t8n+IxjGY0y3NSKQtYsfTBJ6Rbp2mfbdokWGBGRRGd3XYXYVrJI
iMLqXzfJACKBesrNOH04oPyDEBUf39DKqolUiESjBQuMTVjLh3BzTdd47tSgVU7MObPod3U53QFb
zviB/OrM0MotLeNFfa6KPAlCj/anENs7nM3r2k/pIFL5F6JYurh22aYs1C2+FdHnjVfpR8QxHmeh
DTeEqLPELeDaVU5Uvk/mH+Cd9l1Dodu+pXUGEAZ8MytUj8MHY2nf8dfEpsu1SWoM5lTMwK6KKH8u
kJNo0k9QaYMq+V3NRGTsamH+6FqTogezl4a2Y+wJ//CfKmYtLuXx/hJHgdJGKp6tdcOpJQjX4J9l
bHXMDhTJ3eBKDOEVVzT9I/JbSHyLKyZ8vjqXmuPkh6oSUIKN89ovnktwnBvsuiuhi4auLI+9tYe/
5/DQIDi4ueqK5UdrbXkZWrOuedZpxwMzaGqa6zTIEh1mUJ4J3k2tpzPEKBhfGGDJC4oUc1ubiq6P
oUw9wANl1jfPEmmEDqCs+X7X8WlKiiu/R3P6oCWR+nFJ3VNDTqc0IkXjByrN1CZurHiWS37gRkb3
/D+DePURD1R+fyGQVQipc39ro17x4lNLtMEP1vhw7GVzuD1l7q6LVjau81O2WTfXwPatBOuTwGqe
S/LcbSJrtBZ6dMKQmiXaCucVmVDIdmCWYqdrDnfwOqbhY6Vy9ZDLJv+dCrHppl7b+PSzRvzHrR2d
8qG7m/LWvcf863JpcZtLlxEFwW6ZNwpVtrML72j4UVDbYbBAv9pj7QPjQNkEZj4jrtP7mGsr0+q9
VFiKImXzc1f2cNT+irhC+8fmFO4IagP7kR3WBWCJBHE7MQeH/+9aU51690qE4ixT02aznz+DYnnA
eZzRQJaYuboOwGZY4ki+IPyvtEk7Q63zovXBAv6p/E8sV/K/tK/08J23llrg3xjJXOUrRMeXKYaH
0sImanSSEJ+VG3yck8XKFmOicMlBYX7/3vc1uXhD6/J+03RMfCwzv5SS3Gt82/8yqeaLTaB++S6D
TH/mhhwr0lq9+oDqnmEuIvVHRhLGa3qEJ5bFsQCIJdT58hZMYnFpqh3T2EsBlxce+Obqwj6pw3ik
JA116AHL8xUvwtuKsvG02ZBnVdzt5iB+FjoyzMC2Ia4WaA/eXWy9a45MPqs/bUK6FpDO2LlnIthA
7PDfzoq7cZvmrdXQeu0PPBgUWYHXg3mzZRU133ckZSPe1fvrmAxu1pKUhNdrqoVjgTB4K7h/9wnY
DBz5apwUCBini8vf85rT5ZuzItbRNidPdhdBOZIVWjuEtZeZSAQqhSmHKpY7w6W993/85eTtCr8q
VnqVuo5MCSc9yQ7+Akq/M1v7uUoyu99snhMLuDB9RtZAjOQet1z2W2iU0PWTWaF6vZvqXtGYBD3q
YLdAkvu5CmMquWxpGaQX8LnFjcxBLBDTPPxwb0/hesRisREIyi5mYpqxXJYHqA3vFxeM81YgcihA
QBz//mBbUK8IjI6VOHLexUmHOfSbk+As3W6wg4CuG4sA0DF/Z02QvoG111RPRbFDROFKgHWKka7F
rElG9wOh35xxQ0QGYAx6fNoxy5HTSY9cTAOFsdsaBw0k1auAFKhgTHrOkb7G+GF98JLynqUV7oXW
FIr/Nnmf2AKqjLMdoe8vew7MaQkTEIPr2/jC9c1pT7oKslQiLsyW3GiEmc+B03t8rhSm/bTmava2
BdTUkI/aQfDDnrD9voJVspvaFLQBseD8Rm0YB6LgZXMGz2DqSNgUT6Ydy248DfMBV0Be72V/31NQ
+IXajkVkOfQaI0KqV5fGxrX6VIIB1fa8Y+9+hstLXupreZwmLh85IcpSA4B0JRM4epDsDts0Bsej
sDn82260PjOc9DSrv7AG/hiFMnpC6GKYiqbVqY/lJspiyEuT7UOlY1YMsZz4gqG4FzwoOI7xzjOU
E1R+ayTjNO7rA6IUU92nWxr3Q1ptZCLYWEEWCDviXc4Ief/ggEajQpeoThhtl6m18VIXCo/AFKsW
/m5P5+fbNRUxp136WAAV/3QVANA6uhTAyfqrD3DkVlG3q0IfQnOr70zgjF7XOWU+SSK6Hedzy5eB
nucumiJ+/mYy5sKlonB3u+l6qPvLIeQTWgA3BnGcUhJ6nECTfIZ1YJpWhgByJrNN4N5vUaACCUj8
i/km5Ym0bS6WaRwUimEr8Jozvyadw82pMKOGxsOE8GI/WkWfBGmedPNTunor+YXkyTrOpyiFkCD0
gVKFcD+U5cIZ7c7s38VFRkouHmcYB9hC7MthTeKim4JeZ8Md3W8QwRqsG5++uYkp+JXLP3PT2eUG
AD26Cx6A82t6SHnLINoH1wzo/I5GaZr9lz05RqYHFdSGTH1z2tRkwSO5R6j0bzSD7faYEoJP9eV9
/vXm670VJNQxS6xEVwzTYYVMEzu66XWy1zMGzP/wlo9JW32yiy6bIIXJ8mWlW3DXsv3zk1FtzqY4
xFTHMM2E4g3CqwNR7r6uiYrQmXCSssey0hkP4VW67/eo52vzt0N2VPYTJ8PXkFedwnpywoUTmRAZ
34oAJGMee3cfV69RxpjGlZcd+TB6f+bVwMMSszHv8Lv9Wqd0RiLSjTYonLhzvB2+T5nM0VlOZYTZ
QtO4KI/eCcn0tD4RykeNRWfnS2MFv/PSqI/mwu0mFI/CdxcFk0pcXr3AMv7E536LpiyhtDkUAeEn
dBHtPZoiZladvbHAw1JAtMBNJ7OamLZku4s1M/i7JDLBtf5rMw8NfcLTTJFR6EaCN/4sp/mW7Ad4
Rh+ygFpxNM+p6oJDuVRQ9Hb9ylnDm/GhGUzSdjRa5F4/03zjskuLo2p4oiTx/fau6B+U/Z8XITfj
I7WarCPqU23DN7bCtqenH6Me+sESiDbr/iyLYS7YhSWA0H8c+RzLNL7C/IQD1JuKa/SnPkgDP187
ENfzbjtCdSzMIRVqpoApnFCnquKD4hKlSexa2JqTrGloAlkpfyCXrpbwy219Y349CVzcQVaKepbY
kHlLlI8ZZeoI3FUqO3T4Rk1oZ8IhtPpWbHePfDlb4lYJ0LHW6wRpp/ekoINPYN2dPeZveimB9pAl
RB/qfXrzX/NdjfT21nqL33xt4bMWDa0qpp7yVhsWnosCEOMEhOJf77tMv3DUDhAr12wB+jC+bL8U
LQwnl7UD6CZW8xSVHQWqaNQt2bep05itT5QVzaEWXeM8oOOC2uWgLS9PWXS+SKHhSBticSBkQDTn
OehlpG4Z3SYgfZYFmMYk51C7+Yji+Dn9TC41+YAqBSYar80yRZz8t9F90/jQzdvIviECmV8nXzBQ
3ssC0N8wgFj4ryIehvuNvNgozr1vBq9gsMcA0fM8PQL7L6lHd8I1eW6pq6l/kgDQ4i6a4FFmEjmo
a1AGL4cOLLCHnbtHKBMdObLUqdEEDo5ewWhFUQsKcX1JjP09+wInhTFy69BPGVjXh3gAASRKjcCw
/d6pDT7N4H5NTudDFZONtayBB9TBqCEOiUAjDeQA2wRHNfsuHMO+S3E4lnjfkSOz8HlSVJX63OD7
fkhCru1V06LBVNEVov0IFazVxQUQdzupSAACAx2SQQdZeZZUSFouvunsuF5wif1kP4NnZILBs7+9
E58+3JZZPIpeckX1mPAM+CRcaSGlOp0CT9YLVcxyMMeocM5t0KbyJlaIgABQfvhx7sWArUsc9MVs
rqXFkTatlEfM1YHUnFI/vkxarjGFeZysOffLt0ziRxgw3wpSUvDtcdPKIWnvTAeVKaCRJ45zorqp
LOSaNZ2W+1SiBmGSKYEctG75joooHjXVHxwGRR6CrTtz09lmKB6Q91cpV8HgMO1MHkjb88Ke8UVf
sxVR4CCuwXxZR51Phdb+rslQwahWpSmrsMNzcmD4cR3X3bKtTYrD7UKI0okhJZfW0r7HHMdd6kN8
w7s9cD9uslIpj74DWQCPfriIEH+9KnZvqw+z2YXI8t5neZ5s+E/D1ZR+6mkX2rUiVb+QRvuWu0zS
m4+2x7b8KPlpujAE/EJBdPrMkOcY+C1UET7bt7nGgvzOoLfqxIJxlgSiK+uWGiRzz4G+SUrLmt3J
G1uiquJQNLSP3DGa6lyPwoq4+iV+P7MMZ686LkEu1+1krmnhDAKIn78rWqKOLSAbNfd91+0ISqSz
Fq17lypaIBCqqHSPuGPNpsogS7XaUUSoHrgs9xBfHI//WXzS2IwlxohPC4MTVO7M1g9REISGsEeK
E7nGGr3P1LqMTMiK/+dbGvw9SZPRNNayV5PfM/shhNaZBiPeUkbaocD7TNQoov3edbhvnmZ/9bC6
hr/awmkBAoo3fR3Iipsa8JnCZ9vZYV6tViRQADvQ8XL/BhJWQjRdIjRpy4sRuHIy4pBiLrGHQPKu
Ovcwt1VQ5nUhnThLjeXtO+KRVoVuzc9NHj8wphIqXmj8l1YCF3j15YOW3RKv8PycBInyj9aLnrxd
FrD4/vRKDmkDEGsEu7dDA2d3ZP/EpJ86GO5pQZ0nmlEdCmeeb5WcjMR0g/q8tD5mwV275f5uVTL4
p2PU2K/vxSwsHmuunvU9Q/jPcwj/WOm8fFx6AE0RpG3FIq/TBh1q2YFFSEUI8OPBlq/etUUExzSy
Xxm9Ay/uQHJwlIkfjOt7N+PMpMYduyzKnFiEc41RnYlxTQzvB/oGNHXbWasef1BdmluI2Jc4p9f1
+W8Ay/URy9IS2c0LGXrgzZoz/R+a6HQn8Ksu1UTBkO4mz1Z312draqjvwkIhiOiDrFUTqgoFZAod
nb5xoph0F/yddcfKP96Sf626L7KECCfr4KCxzgt8r55r8nkGpdW3RWBnepbrUmm0KbaVVwi8f3/X
RLHnCJHgMqnOdq+vGYtQE0iAQlqMDRmNSR9lp4MbjKKMKgHA8YOanYa8K8mEAcXNUsKnYXXvEaHs
1XYntWHFIbofEIv7wedn6GpuTXUzQw5qT9JVRp3ydK4fdhcZatY3Rk4GDdNYFEyykO7cHpVLMvew
i1uSI3kf2qYZYC5H4AcHeA1mMFQkfg9IsEKbh8Mvlc9zmZvlo2+d41xwBj77BCc2Hh9DJX64J9pt
fD2qMbxNdFquYhOg6h83zTdQWXZjrhLyXYGDGkR7qUvCyM+3SrQddl0pkPaneAQG0J4sHN4tfDeD
HyyCMUCRZ0vfYwEskVzLE2UHFTveCm6l3yolaZpDD+tSmcyd2gcI0XQOvgRdYN6QFE9AVwfIJfNV
7FbuMABya41TolAFE9EG41xjK4hIY0nmGrg+30KrSC0wGo0DypaCmdOTuRO9F2rmUr/6rI8XxFb0
LQq/uMMZmcZ36zTvHaDTscHr0tTjWAJKFl69WRCLi5+ktpiwvY2S5vVFglwOG720xy8hfuP1Yh9h
x5eGJosZtJk7JorbyorxR0EzAUvk/HssK84fYqQbUUiHEcRHV0TkRLoyHmHOPUjyRc5H9XnF4+7N
PB8UQsQpPOkdwqEHBgK/HHBw7AO1+mSh+1CLJaJ1auUZTxAdYqOC3TzfRed0vXBDw0RnCUKY3chx
pnpqRaMGqkXcDxI3Vlku0E9HpTycf8n+fdeYLLE4KZ8EzwGwAd8bPWA0b/2ees8ySyGpGrYYhjUG
Qi15tWgRP+osB/IGq3cWT/kL7CTvHS7yKQ/tV2PBNJrmVjqDdknOFnyekI63HTOARKuRQdUMetap
805H/6aa8Bu3lnaN5EU2Q4SM5at8lfV28PcXhNQdgx41/RCiZ6OvcWKmDH7VGtBrEzOxdKfk8oAA
HR2AOAx3v3yKSSGAFKRYeyQHz8D0bVVd3Fxp3IgRV4jdlYNtWS6NEejT8BZFmp/amR2Fcm+9iqpm
4qWp7F6MapMMjlrtoXP/8bxqvBcuAphL5Ii4gCflnGF90W+lBGhp2QxwrPkVYiI3a6XfNVKqFTKF
t21CV8J09/r8YIvt/diPBSof5FVxmZ0o96guVRTZN1pbqwl9Gbz9vjDK+y/DjcZL2R2HDnY7Z+s4
6hvUT/fSTFZVlUr6XCmmSj6HBS4AzHKrn2YFiRJIw/3TK9abcysAzXwRp+wKSJy2M83Htvji73sB
h+/aAv11zW5ttJ3UelfDGjxZybqDrZHl35PYwru2buzYnIdlIsjL1czfGEF8ANr9dHZqAzO5gpIs
nCKS6q4LfRQGkcAPPsQPVWvlkOwnsi0CDKUVWbY7mc1QgJ685zB4SsPbZOoAdG9hD++xDZ4j8YlQ
351MohQS0BC5EIp4FzOL60bsznRoL2XgIS1qAsuhgju3uDC/22G8kznhDZ3g6m2TigSCjI8eQFIn
XShVOiVKGWFziGzD6L1ZkL3Ww2kUB4XFTxqeaJvpQVkVxgvMEG4ANPAA49sGIHXVMpspRoj8iyH/
wZjfqYuhuERt79jHkaZiGH7MIVI8oBhk8zA1PVcLFWTuOF+BjYzXo5BYTxrogQ/tSBM9FZqYGrj3
4BA8SUa+mBXdYtm2ZNhc7VTe+3cH74fAS9oxSPeofG7alXv/ZEjPJoiEkaxVb9xmw8S1mDFOS/o9
5zfZY6XuHapQx5PV8/fJBkYGKRWblI4X3xpB4lp6SM2mx5NbciAMQlbEJntYCutCIuxHcEKaNu8Q
pwyKoik3g8rxqtge34pjZpeSR7Yf99Ba41d0LJT+Q2+3eASPQPMXf05DtN3MejVSDoCOa0PVZcgs
e2nFJWbDmvSFmtthK/exvU7lkQRUwyv6iFrmIS+dj97c3/4Jp6diJT6rnaHVZVBazcaFmobgvrbl
EMbTydXatRoo0pLUzcot00+T+R1CZA1k9KioQ45ryCKRrOJDzzlyoi0LsiZj0Z66stov453hx305
0Qf6sIzLmzOWdxUqTMmDVHrHdEMQBCoWUZbnmJqriez7GzTKwB9G57ihLKrvrOt9xUVAnx6Qf3/G
LiJoFX7VGHeIX/AEICt7QTU8UMh6+fFJHm/NJcqZi0vooAf0ljdDkmvNBMOVLA8VdzUHa2DdL2Pz
PPJp2bowmKbGldBNwiG/LRtTr5QtI+bnE5dMc0/pZtWrYTZwCAt+OtLlnsoscpT7pPRcursdg6mL
fjzBBvxiBHgax7Mo2GFJsX4gq/fmc8D5hvN0dsUxDx+bFWfIczIOK0+VJWi9s93q0FakSDP4gG6S
aWSX26LveOjHhA0ZN3nBtjlwHTHeF2tkP1V3Rrhz3mpWNyIu/ybq5OcWHxOi3edb/ANXosNQVm1D
qQI2qdJgrQ/D6Q2vPlIake2sBb6uYCeTp0JudW+sPpv4xGWcYnhFpI14LFlns6VL4p78sxGZRsHR
pO/kEEGLKClOao4a4dYprrhtyahTOKswsmlaEeEBcCCLeBvX7JuDvmOl7DhEST/yS6WjfMrS8dX3
xB0rjHgEBPrfDOAzSJRYhQ2z33iXRMyfArWqT1rj7FBYUiomQDVjSRodaPC8G+wBsLO5CGMNkmO8
Ff6xhEClRjzREg6Dv0sbYW31vYjUJU7kh3LeDrJ/jil53WdUHPqeo1nQO823skGdKImI6CkGe5HJ
8QcAZKd7Mhf8zfcEhcokDOP45HuEpEYyGN8RXej/xTM+Lp2A0RgC957xHaYBkhRhyoAhDTETLzBw
6MoATMP9MUWwFq+kM+oq8i9ozqnenwxowTJhBGST5JunTKt9QkXEzWe6w+YBsTOHhAJO/Js+W5uE
w7OG9nuhZpe1vYLra2k6ISesxmHwU4N6W76TQfuklgYS3Y40gcPyfJvfJnFnAj6A/XcyvA335pRH
nsU0Y/y29/seKScr9pX5w8jkuWy26jo9EOw/PTZ/XBWHhr2eBk1OsC2j9w1ooL/1ndLZWrNiFlR8
uTwCBFdMgeFGJgKoFbc6m6q0f6zCsFl6Wp8DaAzyuBs4yEwV9FzZxB6nt6cQpVWkolz/rNRYTaIe
oqlwbeepvYg32n30AOafHoUgRVyJIZ9afTMuYt0PeM1rHhbe5kE8U1y2ypRpZ8ruZ/aUpI7BLVIF
GYLZ1z/naUN+7GxXcSgwGGsfLrhzpZ68II80wJ1j2H/WUwARRWZjsRVZV0yaWdlINjjv7NICWubc
9q1j9MK6f1T+fV7Jpl4CTC5uzpObI/Q8XokvXy3NhjYvAsKslR5hvzOadB6gYYSXGf4RAx4+AqR6
884aMfBxBbdr1vDPESBErtidJgG2A/5KzRfoJcLL6sZ1i2rXn35zJtKo70bIwvUmral6Uej4Yci9
p8ixbHszGTe2Tokv0fIzIkdxFRt+UcfQCmRetaCVQas0BHgkUMxomyjvkooWdKO3q2bZnB58qHvz
zNeZ95J6FZfdR/Z/3zeJyalBSFeF1/Aj0NUpyxrNhGnJxNERPEiPerIHKIxS7jm4wahvjnzQVTt2
1IMoQp3D56YnSc6sr531rawXHLTlRTM57uo5BoIWiqfyZv3HlUMBeZFVM30zlUMlSRH2X0H7i6Yu
ZjQR5brBz3mLkZqdI4LjLv2JRSQy2g7K0oJ/p4k7AFbDQRVj9Olz9WaxZf3tJcxIW1HccQLdagb9
WGNHMNrf877z1WVmSOkGh0XBPDzf+OBKe13o0EiAupVuWnct8AcfuP5BbIfZEbMW5XwPBUR1ATJK
IRaW4cxW5YpuXSSwyQU56SNi+cuV35uqlQyHfhu6oRHBKGMdiNkglBoOHViO4osCU0Gx19HOda1c
qhW4GuAl8h8XtNIegzefFRLhzMt0Antg4cdxiyWUbs9jb8N7biVZJfNwMCmrAih2vm1rybJ4h0yV
kY4sHt8QCQx6nqrAiHhP0noadtATZYGpk2Pf6YD8zFE8WHNWiS/Oj8H+SWAyItpyoMhorxmJ1zmR
NyF8LLQCaeZmFTACR9b130o1YVWIs1F7ohT5vYyUH4nXM2c6m1QHNlVONjDZfmViiQ6XoCKfK6Oi
2z4faozy9pJoWxtySdF+JM/tVLp/c4nxJ4ZmSihX+tNfjrLRUALOhZEEudBANjK/ZPnNSju5BdX7
Kp3dNLA1M/JPDN1YNrgaLk96ZTDST68h4xaW1IH/e6Ee1jRWkby63XvvkdItfIvYWo3Axv0sbguQ
hY3rwPZyeGIUtHA/Ma9A2wqejljhTtL0rwj0eCYWs31KfnP2kqFva3ixne5po7YUyox39lia5lrK
DdWuU84KgSyiHrfKJVm3sQ/RtXCulXvQdIfWPdqEBoMMO6LBEQdd2s2RSCL4ruE/2RLQXygNN/Qo
CpqsZqOFEp6Ohg8mV13EtyoypUA1aRH874F1BsMTa6ccGXpMIuWUEwSLrM50WocXxsM5hvBl2TQ8
Qsh0rXPVw38WD9HepEn0WhDB4PF9rhCc7oL3uR9EJKjpJQICaRl5BiLqmFErHOl78t5hfs4Yi7m4
vCQBO5/zOU3QNFl35PkLWvDDP6AhZFaISeU5Z4fMyQQo3cO6BOIo2vgLgpfk2N1mD7d0WfJZK9lR
UvINa3dtm68ZASEDLkwrsyoYSDgFzXVbrgtX7T3SDt10TdzjCKANiFZe+UPM18UGvTT6PGI1l0gy
+oIOSRj1cdUEAYTun8D3rmO0omcBiz9mJXv+FsnHR2jy0K5rT1STtg4a92mp+hqW/0o15SHJBfCr
ys28Gzt793cw2wI23V04vxaIFRovF5wIdXrt+aHYELshDVFMsWU4P56SsF8fpt/c8qehIQn4x2Qv
4xLNahGvP93kgLqIqb+aJushiitKH6zQimMEiloTe+R3uUzt5oxDHKIsCYsJOsE4/bsdZuLVdntq
qHODj/PiXHLxZuk9iWxfYdQpZ+AEIUM5VkSn6SpL1FGkQtu0jXMUAoxkgWf7sNi7cqGuQVIKxQAJ
nDirm3Hp4d7+8V3HSCwzk1eaFUDst6PTQMwgHdGuxo+aH3xNdS/Nru8JR1VkfieHUmmls+slZBOU
7E6Bl7ng+G0UbmjFzN8TqfZZp1uZHMYQYqfWMjNj6rpmceRzlbfc7jl0MvK0eWRFQqk6Nlajp5CS
q+d+xgUDOVUDHLCULdmHox7DwJNBJNwMCH29iFrbS77xUh3p9agQX85X6VTWkwSdpUQy8xrssEew
flJrml3c40tXowr27Ftbvlr6oh2M7Wed0unE3n/LgqvFee+tfO41ZrzNPlEJzcqG7R8S7oKHdCXk
9qvJ9KypqJinNxP49/ZLT9M3+44OcyWJ6TWyh7Vo6ph3a8nfyVtYm1cano83IBp6Ab22kwv/2zXP
hDRAI7RZ5PXISnKR+T8HAr6VlQJ4Ng5ZRu1RTVSe6e8XM9/yZXJgwyshLrpHIGAo/qyI6CT4jEyM
hGrWOCu5Q4+uipfu7mJOZGgsCAeZOEUuCy/aiDOgO8VgRzREBplJJKR0kB4b7YJ/vA+EAShDu0dv
e929+VYLtYqgBoeETJVkqvuKTu/X2lrORzDCW/tL4WtUfLHF6f1Qxc7FBWaOS+5Ss6yoAwFO2DUh
mzRDh6KHNwF9LVvnNEBDECCGDhCCtoJXrdfHN1UekgOATp+9BRaV9cd/mSTed7PzkCW3ddVp0UQO
j8I8RwE3Io6Ui0LoQrb9rlfa72St3Bjvefh6kI1MrA6YGd6PwAXMoNGN1oBBjaGDY/x+ErSEy24l
SsrsoCRWX0I7B79dVxjjHIYKcFrHT17nRO/ZWSEFay5BS8qh7ctVVg6qjkiWz2fL33yrW/z6OsPR
xCXL3tFDoffrPPDa6+XT1yGyPOuCu0XFv0n3OFMcE+Z8Ujj8oMb9y/qtFmFPLVcMtPVyUyiWAPQ4
IUFPjqFFpbxZqMfXUQj31xkC/mN1SyUxih45hNMX5IeAedqdn3a56NzU/rEZp1brfgR2FPD8ytX0
oiWyq6+NXkxQt9O26ayI/Ug9LcSnpikK0L8YhO/9jlfD8Kw/erb86MpRz+FfMsM50WwI4E7iZfXO
H+BkykwBLX4Nvd6aTYgCwtKcj4rYazOghf/kxle7iQ9Ze6kDCUr2UkPACeKdGkNF5pytyonn2izu
eQ1sxxMmKYqMjx6IAqCnXVLqFTyN5boqZvbexvMgbCS2IuXBnU/TuWykkzQXOVdUj+Yz3vbj5U2t
MEfewNzWP6T2D4te0UlpvJ3WyKg+sxXAmK46eWtKyr5eZKLvZHulz9nJb47LcfUzHfzJyLtlSDvk
a7NjDBCicjI2ttSei6MVAqEA6C5X5p1ftcq+TeESafQUMtgTp2KrVDOStca50KvOLaeXsIjaZtG7
CXcSvkKZ21auX2obr9cPYBnJMTuviil5ixxP73KjGTr5Pz0TkAcSR6jqZbrMoKAXexhHlr8NPFnn
yzo0/eAg222H/eyrT9AA9j3DlGa36rD5Ulh4GINSBTaiwvRfsojOg7HWQj2DK7oWj0lXRyYYnn5Y
9fh8beCALJx2K404cqjS4x1OYC/ZKV4cokGY6jBexu9pQHKjSttTz2yj93hSdCNETM6VBy1Kza2M
CX03tSgJ7a54uPj/Atum1JXhcNSUC6c8PCuFXGbsV+2/Ze/A9njQfDcajFQciEWQ9B6jrx40iEgi
t8tX9SisfDS2oNCFCLmjTUvkJuEvK9uddwFerFEo0FnU4Z53eHA/ASDXwhRGTkifQ4iTlcSYnvqo
Rshxai+kzXVzF2Tvyd69U1vVHpbcfFxx7uQ+khnG+87wEP6/ULALyF1NtX0PbU8yc8zX3OGOhDmw
RkDk1uETyg6mKleUdZl0adhIjyLW2QNTxokes/+GV5hsOOzn9Inv8jcw5fG2vL+1AjQBorWjcLUz
TjVSNbBLp8WLHNaX21ZUeI15KHOKmNDSbhE4EftW+qe2rGthUEVlWoWT3E4f4K98rpZO2W/tp9Yv
NuZOvD/LhzjHYzxe3vjSMSZyiVz4Z1TYQw0T7PK0JsOTJl5OioFQw2WdO+j+oml5YIaDMYhkuAf1
LDtBEa8r+X3yBC4rPlJVsHtcE9Pd2J4VTqMQNurd7eYEumMF4WN1OuT/H9brYZtayOHcgA2ap2Oa
Lxfv0cCtk8F0Z36FSb/E4gLcjRHymBtrZYftuRtgwhrE9g7AiOLSVD9vmZ5mtDNIF+bsFhG0sLMp
a0xZxDDO5pcjwJllbfUSpwkjsPYcfb5RGXJ4Ef7b2mSmTqHGnpZN1zss3aURqKRfhThe3HXtFFjn
cE9jarzNrxtT6i63uHzd99dxNSxTkTMHI9qSMzdDfUElENIz6L3aFiGtWOrYGAm/YVMOyPB6b3dy
7FhTUjh4b/hwkGviS2PfYR1/vQaCrmU33mglm0pKQRkbzlmH6twNHuAdkWfq4jv4HlwDEDq9D75P
MBQ2e0Y4eIVLwsBX4ULeNYyX5QfsWmlrH+wgK/5Bn24rmhEnKkvhYdSw4qnJYi7Lu+Wk6SRup16d
5n9Em9UH/F+CMZDzGaGIORuNDepWk1ZBSo7IzeuK2Xm4JAs99Fwyer6BrDeeHtDWUPFcVNHyHip/
sfygxeDqW+yNlt73aXMFTf8cYzlLJxsqJjb8lgBHvHq+rEO/vIX5BW4dg7Deaut20pz0kfjXMes/
ApsJEFfF8e3z86+9o9h7vIbmGPiYUDT3fp60eS91IPAv34G4HEZo4cFQSjcO7rGMvd7NFS7MdPfJ
aBTPBcwIS/XGkw8iJWDhEn03/ksSmou1HP1dQ9nwAKCAk7y3UH4SUSar6XpL2oSWHkZfkNaXw783
L90/AaYraIyCGt4aAwc2yMv/BFMgrgOPsCgdlSm/ZXe+S29oa6FvTnapiCFrW5udwjaw/o0BH8qb
QAMGNITtGoiyen2ngOoBDz4UfvbAOhTjigrwW43Qn7nBmL2Z9lHrhCT/6QUydcB7ivKLln+DfeKc
incp2wp61TOhRUMVcvd0k8lkLerpUCYbuAs+TSL99JLiCpKP6JqD2BnNIzEhu/MXreQHB1DbSd4m
CVI9xyBBfsMCj7X4elXLUBCiWy89GInoPavHpUWtAW3rSwMkTbYXxUmGOpNA9PN03uO2Z5aI22Od
kkh11v4U2bXqAS/G00J1xQjnaRel4/ScR/r6RtJo6pDfLlb1EtzEq80dTpPJqV5Hr3kB2WkUHaoD
jfrfEE/Ziqm1kWBO1qKN5h5YmGC0CNYF5Cg346bwljkuTRHKPbHpHLWnA1Sne+PYzRSj2/tgTf2N
pNv/zoc/7q6Q6o/EI2l73lPzFpLPUp2WC/xFm4j/X9m5Yk/yNg7KMJFk+TzA4qJkmZVwyWM9r1pN
UNeV3Kcwu/vi4kZE/hiaCY2mafOZ/jMX3KwIft3dKPV69wZHWtNLMA+4HobIZ0GIU9c3LliXLWMM
F4P6rN3H5lPmxtnqDpRwIvxjtaUzikzVXtMGQnFqzXp10tnTXcYocKek+qF4z7D3+qIoEp785DGB
NmXk9GGrHPtiJymEGnbNxcpLOMjda6YC+sB06eWQxcf/bg83lla/eZM3SAu0B9cJnMucL3zUWgYc
QNLV5GuIZLl6cq5kO5+iluHXCHe+utXQbt2TPAFeYTwaqj7+vZZvy9AE7wLLEZShFtwS4za3uFpO
U5/s1KWF5PsPY4BVsTPmv8JQKwZzyewdwyWTLhVSBrh6qYeYTBoQZxz5wKXlak5LcVU53sVLcdTA
yM471VD1++/dwyjTN8d+kPtAnn4vIe0mnr9v3cT8H/2yeFBR7pZNMXFdjDVppDX9ofbmy5HSVklV
UqMpjHRoPNVMBHl6YB7w/SJI4uvlyLtFzEkvqwM/aXruX4JF7IbArJUx/Hp1QQYc4W5w/py6oFJv
+G/LJotd/sVq422OSO3GUE31BWDPX7I4Ejgc2W08bDXXIM2DQYHDF0v/xhnQW8bqWN7IEy9t1GBY
Khzp/9wQprFM5r1eg94CEXteAYo8oY0/AGU6gMGNZ4L0Qei0jmu1p7mrdkCS7fJiuoA6y3DgmSzF
9sBIud8IgpPHjFRgnz4RocRP8lU7otpqkjn74W1lt82Z0U0p/x0Ex5nS9W1BbPANhsnfon+tlqW5
UGlgY6wS41VtyKj358A/mvpcNjdg21GsdBW+u+jkB7mzqt9Rms1iEAXOvvtgYr5zmi5dNSFYdjlw
MEZcTTZdiJGIb+kA4SPJox2qg3IMepikUTF1cxOklR3l1ifoyio4PZ7/acbGK53recB9Ejxiu4hb
JYVH2giPD3j4WirwMslFn8cqcsFBoqlp38tf5Cjb1pKByVpJpW1KzllM9arvRVlDY2VZbnDQQ92M
zFCI4w4jssTUjahegDobzwFql1VyTugUIm0HcnvxG/eJxvi0/thEUUwLJRNu/zzZFWCO/1BiUm52
ExEjegqsog3dvyD4vqqcoxXqk5dMGe9KXJkKXEcZfqxdDsPBTLjp7961RHucjbt8fO9UT6mtTbdw
Lwh2NpbEZhABDTfelEvLHm61T26wk/U/HBsBHDnvQiHw1iNtGk9kDblay0jDPTmadTQWP6i8hKnI
wSFGMQELCjNdg4GxBb8lcqRiTOJKx2zGW+fFk7mCv0ZXPwbrMamwS03SxDwjtr4JjixxPSup8ORD
hPksKL578ukkiru90xi0Ms6RTkmuZqDxm7hvvv0aDThDydMM1IpzrqbO+J4nymfdmy5nGCtDPWzU
cl+gdOePzQJCbZs9Fe+IsLwC75ObOacxYND7CtewdDekzRlsO5iw2aQ3b/IJmjGNkTlOfmO5v94I
nlWFTuJuYpQz3hdW4+eD56nrwTzPRv+nVgAMv8ifj98izaU6Ym6kgkd1W8ybSA3ip2IPxeZeSOcj
ojlJRkVBI1sbOPWam6kJmNr7FUfKPD4aciv62TFO9Hxn6s265k74AMSwRRGU2hkBx/aMsI57E0pG
q32ZF9wo44EtRjNp0H38YXf3u9h4Vr024vrt/X7LvaP2m9nIgYFVJI1CTCdhyubiQUEjDvPML4b7
SXyHpgKFTYv1tk38LfCbaIodRPbcBwWqWRL71/pGG8qEZWtxvv8PaJMINAgp1Z1iSN+lGTu6tG8t
4AKMVXoUwI5RYQQ8BV+syCGXCQhG5dynPSK73sapfDpUUPngrui8bHple7U+BHRG36L5Zo3v2tpM
KUpELKVuJpeXDBrPLlSxvSWb+ZVBRSs8+h3RvD0sI4Sq7ClkuQUS+bHztUGdUzOeNZvqoLx52FWG
6PM03Gb+KDz7VkvFXF+/bXdDjHchTotJDSJSd7WhK5Wqeq9O6BeeGlsEg/VQ5+vnIj6Ybk7QZy5w
1NK4rEXgbrMHOJCtYmbwe60bSaOAD+kcjXQNpVj0FtBgxPkuqhX5Oaakc3j+KUrKLB3m4IUAkO98
GEHVGXtTWnZZJAeYzUF1TsKm31DIR86E/vdhD7EoHbp1pLo13f/vNj/H80SV96KFCgYGW64EoAli
Qjf0MzJURZ/wvZKuNo4M6nXRsMQTO15Kr8MTFmBdBOMqvAFGV0URqFtcjZiFecKsOUHV9hh4vUbL
zUK9ka4iySQE8WUb9Hg0DCasYvwTJDgMCMuT/Xzu7TZ+JTKgeN20GYB+TktpcewTfXkkK0okjyKh
M8+Hilf7ItO4p9MljRlnlDXBqhGSHdC8PqNs03n46RjkyJI6PuJtmOu2gx6KS1TytL/2zlzHSWWL
XFQIw4lksSJSJfY5/O5n8UeUwkRSdlWMlmwjf/g+fKA8AX0PDG0Yc96dGhgTDBLVKMJ/RllCg0TP
9EM0rqC4N9H9+ORC4xNZo/TeiW9JLuh4ie9KUQs5ayBPFn6/RlSojcjLQRjEq5Dr5MEl9L8aml+o
BGejpjTIalqqr1I7ccMGL2cRhnA6a6mt5/cHbFMrsJ+q6v/xJCPyf5VMzBSmCC/wEw9dri8McmY4
HDuYrRMGVN+PX0oKNJjp9U09TMkmYDi3/UZRsSUK+xIPcTJEM26x1nLeRFQDOYmpMFuLFEmiLpL+
4g7F23IQTfASdZ1ZW4agoxLWxCa6RKig2X8B/JcGw5Tq4RUALsnyJ0iMWTSrkfnW4fccXGTmmidP
fvzL7UbCCsTNOq708X4Bc2fEb33Nwk2HSvj37kcDxQTLx77iZGTsH5KdHfrvOlqgPynnjXHRBJEP
XxAIR4z6NvWp+iuAI0s+N/PdKNWYoHXryaySH3G3unhLYclt9tCs1mVo4mdbnPVplBmNnkabQJ+z
hL1r+v6q+Do/AD+8iHy+VhuLd08k0wqboVK+/ZIxolevHBzR5YsUAAvZ33bILT/+p0OFS245X4Z8
hD6sUttaMsErS7Q5x9QcnRc5Xb5QqTiavjAgebsw8trSsvH+myqEHZ9+4XcH91QOybdsjHrQ6zSk
Ko+Jk07AYV1RoELjeEQc3sZGVAh1S7n6e35iiINAOWPwu32DSE95oanlFOukTegh9azgCf7a9q57
jc9kRQ4U6nnwWRuvOvQdd3go2pwv9YyEldnemJ+GSHk4m2qoD53lMDpyx5SyXqoDF0miM4JfXMzD
m0gwkS0f2mYuF0ptDeOfVO6l5XoEeZy5NP8P8zJUdgniuH1dVvuZt9RXgixPZcNLiYGKj2OIYq6t
n2ZUb0bnxRFuKUzVRRP7qtcW8NZC0cdZX96xvAEpjkitflZ5GAg8iNGAUKw+Y3fdSSPTwRvOVVej
yRVFjwa3bOmDX5UJhKtQrP1xBkbHY3Ky1z42OY6vlrpmZJsLvOJI9TFF7YoP0thvCT34PhahUqOm
Ey1BCrWdNj+/gucf9nIost42F688mtMrjEnigjj/c5Xqbfp1KpYKSh83sgOvlhe1STccDNn2YIRh
1/8TeSXmpsXx0h6dnfZBDWnuCNSBybT1crjIwMNEdgKdstXXKff7WqI9E9sksSt4zFClphT21Jm0
fh8Z7Fl0hHFR4z/hjb5tksIPPMbcfpf0yX6kvJt5nDeQzWKXVFPz/BAuS57Z45xfD45arWSb/FBL
/l9xlw7IcmX+DoWsfbpuLlObHQvtrus8vO0QiSqrC+a0/CMNj/SdIAfMdj2FLyRs6ckg4MP+HVLa
ultkaWS7EizMAzj7Zp3pWY06ZGVpysYj/FmpcmnSaclyjlC4/4MoTx6wkMHna4FFfgdEKZF+L9rK
8fx9krlUYOzBy/vB9IEMCSK0sYDXx8yhwXZZQ1+f2PjunTKU7//hqQweb545qwtCz7vVXiT5z1W7
Qmg6rxjqKSfg1ZH7PPkWeVi1YHQfSz/nOpWLbsA2vN2+zlHN2WBzKkEjwRNGlY3IORIyCCvvezdq
RcRYzTcPqI81u3MtS+73vL206JUEXQLSRgq0XaOG4cmzBsxWIrryqddwl65eBzFTozO//OoSkt5C
6IlH8jdQd/OepDHRknJY9B1otDiXyWnKWYs4LBWk+NFkRyE7qmqwXwS8Q6HsO0hY/vGQd5Z0yDi6
fq7m/lvpTPyS65XJW9lnQmMBHRt7jBCFANwtsy9p5n39us3Tc9b14L6VP1xnRsRNJ7HOds87CV0X
c72gt+aqwWLDV5P+UY+fbChl1GnMNmWaAAaKa/KwbXVqypVpYZCJuPvXwk7yS+HXvzroNH5DC/4K
VZqKsYvbTQoIB3Ib2ruWZpfD/JdqXcc3exgxvtVUPurZMLRRtRQHM8o8f2fyy7qmwyZV7Mo+vfxX
7DDVu/zYTMOvYjztTrUrMiA28HPK3yry6J8/MJtDuV/wHfrqL1Nzg9WHux7CYzZLsEWTi6jABxW2
e1ORnex93IL4hd3oBTCJs7M2Whu1h/aq88UR0jnVgiDVjq2ZM384PoLzSd3gyNZQNoKT8Wfp6g8d
ykOSF/7Mt7JeL27ys2/fLsGqSrFe9ewQdMf+j6RCQ4p+n+Y3BlgV7tSwozHPOwqofRMJfwR/F90G
sLM42Rrw759aGZNpnrA/GH1zG1p8+d0SEV7uk17Vtg5nBk91ltxv8ENxUieR2xq/LmhEpYY/nh8+
j0MnN/25hyCxXLDSgB1z5P8UTURUE9xpiD9Qf/bh/uIKLnf04u5oFxAaXmWgF0iqxWeZue1QMQu5
Ya9iT0U6nYA0trTjrTOakCH7tWPqMfjGKLxtovnafWy8YlQLUaHWFbah09TX48DrATBhYNYSHMCh
jWhnhczEUjb9JTEAG6lVvMunMbi3dCHiPYPjWiiFl6FsU2iRz0YaIfXbenkHwJwGktXB21R6RZcw
qozqMvvgJF+D3kpok2hYLjQikgzrLbIfGTrUE8nV3ewCbaYzYcvzS0WBgt0bvXurj4OKXu3681Dj
A1ja/IUOn5AoiWfl862AoImUB0zvvlMa9/Cj1J4eqltEl084A2ZUZF2ul7VcJy1Q9B59aFiSl20b
XHrRec4QGAByC6e84hki7lUPnuBZKjGuOVnhjTYfZyaSd4JlUV7TZd+C0wIb771flnd3Y1eKvBq3
bV2A4zFjC8vH/RQPfVOrknlsGLXnYIjtC1NCqMDRjQHjbpdbZKrpe3IcZaE4hmBZUizKQY5JB502
oflaFpE31HGTOJOPyLI1EvvXnWe2+kQB7AeZ33+/ZlU0DY4DZp+7Aa3i/fy2HZ5gHwJoMsockU8h
6lBbj1HLuDlq4mQVXtnf9dy7NaiI7QkCaub324swBZyM6ooM+DgcfnIaXlH9TfvBDomARoOhBBiJ
ImwiCO4SWN+xnUKPVMH3DAYzD2DzaxCMuQv2Bs3KIlOetGQn+uaTKsIG4liYqyKnDKXJ41yXS3R7
xGhMe0/k8WxyUVIhFEEpyMNoEPg2hXYnj0+JlzdnRGFJ8Bz0igrpj0FSXcmzwAeR2J+tMQWpJVrf
Px2HzSRFujX2s+joRMniNBYfmyjJfqdhk1zc3t/2tKI3ue+gYuNiELF8Q/SJsb6MUSHXH29qhARS
Ej+RedFyb3g9UvILEJbhoa50dsSVCmLKySuQfjHcwcXZQZC4g3VhNieSIwKq7/wldwenmTmwQDfQ
1597JuiashtOAffU0spPUwF1HPcfsJR6mfpggGcBKBt2LGDmAwPTs/m6gkw3qlnZkRjrGjNhnapf
8xfG5bsKS1z9FpNLOIuJvGg+KvJHS9z8QHXTBT97rktAkQN+JAIx/P7qmiBC/BQPDgvvBlMwb8Gg
f3JGpzk0SIRBnE2AUBAmWVZgh6UK+ufq25qtvDNfxdJvw+Kb+6VxHB0Xs/UBBelKEJxTcbX3DYQq
7Lh8vtvLYxReId5zkS8MknsHMa2RHaIhJkL+4PIHDebOk7y4WcTni4CmmPCBLEx5RFTkBaSYB7iu
4EAVe9vDCpQCi+QvpG+66NXBhjUkOO7mx8TJzondRFSFB78X/YWk6IwOYR3FJ1d5HvxR7Emmmj/6
CogVhpJ9aPu0lZNpFw6UCp3JiPmH64PhEOTcuOCuJdG62LLMCTWd6dVMH6RpYHdKrb3IBdsMfnxA
HZIGesuqIoVmvQ7qjNK/4dj/GoFBTUFQ4Ck1W6UYxOaLaFNlDDA5zxwwgk0cteR5VRwA0jPU3LjU
/0JQGMFJTDjijF46TjjQn+beXzmTm6DLxXxh42j2WqyaFbj6oyBJwbKSuQvNbo42x/2OrACSxHGc
AW+PUlg8QxZeCpmQ+mdP1mpdhHwzay/razlP0up/zu1ylqgxwrrFeOYct5tdAskZRTRmC48Eov+i
W3NOISQyZf6sqiEmeN9t9wfoKKTaVyusZKRcZQNjxfgp5Vcvn2RVamuMpQO7vT1HBTfA9SUujPyI
M0Yaa08u0hNa3zvJiwxwIKQEfPD0nLLU6UNEg6Cx9Tu53rglOqnc46xuji5/PRjAOT1VtTKLJhgI
zfRdD5BNRf+DroUQ9UJpaMuea+2sqKcoB47YyPa1Dwyb49fjf2WJ7UxRhKAGXEX8xgakrGPhIZ4i
n8XjBF9kPku2mLH/ypVOg/jgMyjNDtp4GDNiDA49axM/OZvtNqL2qHTBEtoHqLQwYpV//sEgoSFC
21Uar41XDmc49wRm+HeszZhHhqAFi6v98XS2m3j7yxjhWPukXn783SkhEV38iOpJ6tiEXM8C9BWu
zS4sKuRknBJYJQPpQe5i4hWSgLgDRHAwbWYRh+p3eTQSFngtraYRCgZyi0pMrRVfOlXJklKHBxBA
guNMnu5up/zSsYzHONq2ajqDqQgsqvpAIjkxXOWT3oITEw3NLcm2qLyBdS9ytFxmJ3gDU+Wtoi/e
Ud3LBHFDnmFoRSJXUIvqD5zWIULWQIgq+N4mfhKzDJfHYCKBUGUeZD8OMDTpz16kInKzbviXPXE+
gyGMeDZQV3yayjjq/Trjr65InX4vOOOyV8rvEUg6Zd7Sp7oAn1unvFQdllqPUvuDFrfl3QlMmWF6
DVpovYwLlcD6ut2VxBYMSygbfmYCmzGH+Y/FD3AwbL0jy4Fjs9S6WsjRLYdEm5GCgqVLYVZwpqBp
qXeP45wVvkjATMugyTtHQgmlP4cbnnsEehwRRcN2DCmo/rWrC7CO3mkQtv8xi/vTzgWbtIS8ZOes
+7ROM6X70P6BV0ZSpo9WKSzWSjRi0tZzTXPxqxRm9bTg+/RmKbPP3uP0MAjDndC4n+F9+0oMqkpi
phUKesWiTnocrHznhNBs9kb9l2796ybsXWurJLOQQo5M/8nf5kbn4y3W4ZOP8HC8JtQ8ND2T9bXd
x4bm9hUwYG5drE5rqlbntvqnlCNakRssohwn0SPwep9Uf0Y1p23qoxYztaQMEBd0URBi56+wB1W1
GeIc+iKYH4evVDAa0jXCUKwJjsitpPzcgnEU+HPlZUQP3Sa+IGkpQZyCiGShkDwg/VGF9dBVn3UH
hyV5hMkZGkLchD7R4n420SaSDlMPrk3MvqjiFeW/EcO2h2rhq0LgqNMP3jXMXykDBmwPs6iIBiQd
Yjwu+wuki83mZGnGtzPkkrNXh900NkUnOibCWJopt/X4Fb1FRFeWSFaF+nViNB56G2Zyq7UexiwX
SgHxE99eFPpjQe2rdnxyBU10d7EIeP7K17jIu9Q+thiZ2ns/h4VuyNAPNGCEn6R/KngDglpGlT30
nQjoboUVrtQ+3JVp9edB3mdOlg7BBuN/onE4FUeD5cK6JBa6obVzuvngbX52c3JxJFxKZBoJRAl/
QtiPcIEB8pRTWHXynY9Tmky0iyTnUGAuxs1iEPlUEfFO1293gvbLE76RH4KxyU4rI2LmiuadN9gx
HLj4FKzgU+QsgwQl1Spiwy7APTzUhZH2tILXQcUIO0hHpC/qxDoNSG8AGF5hAK/Ed4Rwcbsx8+WC
9gMSQOBQJJJlblqS4g6powO9wDurVYUH7uX24u5yi2zo3kQIipdUAjfjFLx+HprEY9QMSQpWaBpk
c4pK+4Fk9R86adpE2rHPM8O8hRV3VSwfng97F+K19yWVGIxHt/C3uSH01Uol7bNsu65S+coHEfeU
CKHchRFHmCPfUzIDLltgH4ZFPNV7AQi/INXyhno/zu/VExB1HhIRZJFjUP9ERRUgWn+/Y7SS2xgE
3JIEMo63JL1FPhDiIz/w5YwPz7cdDGUsfiOrwnWR36iZbtBp0RhXWHsqXk3ohEpkGwRhZHYE89dc
WYjKuSt85up8IuiuXgvZTWarSzSL1+QaaV5YHW09JEfkXWOP7C2UhPycLPvEFTQHre9bQmJGADRI
Vos12jlzwmehryeZZa0QihgOsuP0hxuyU0cY71EPRRMLW4TEEPFdVggi9gelmwcgMlZPbBehxQAR
MM4WJFg55VHaUb2M1jvdEyWGeR/6bWAaVszAYuPgxbAaoXiTtRxVrGz9Ooh5uvdBbIaKYWczD532
QGxZBUZlaMcftEzzEWWuRZbKxpfp5mu0QfishrN3rB+ddfbBtrzYJmXSwrAX9kNAki79QrfNfDxv
q7spXV4dVs6/ESHN37z77Z9XjW+YJZonawq+2fuby7O8Uce/t7kwewbpQ45+H55yJGsrk9XkSoda
6Asq0JI0fEbm9RwitQPysHtKnrEUlHcpbZGjg+2z23viENUZKPJRmjcup3Pu0NZ7qr4sl2x532HC
gx23eka/IQRtYob1gYfGjg7rsRBZ4L7EVJLH52EEIo3a2okAozd0ij9xfiFRjfOAnXWLXBa7iiZn
r7+r5m2X8lOms2HtYpXie8frP1GFluhGVzU6KxuNok8BYRvxfe/jN2O1EpgfAmBdarn8eORWt1eR
GyZS+7Q4Q9ndm/mvMtTcnw2TNfTR8ZCjhj/KkrU67vhPodLIv67Rva0p9dnKSL+CNsTkr2DadpEa
AyAAXlttgnjuZLDoEhlFDLbjFheROPz4uC1Lndkj3gEE7kU9+DU3U/68xqaotjCCZ+KPx75Gam02
8GbxbScDnW4n+KjnPJzscII1lOEu7zvnw1m+3hA1bq/FR1y3EZ+FJmmGNHLcMSetos646UuzLm1Y
GSRdkXZmsEenLkwQh5xQBTGKT1db1HGiuKVLl2aYBukfn1iyUOPnAUhm1sCrjpfXDV2HbaEJSmGY
QK9Rf3W/Z869iXZSDT/VuoEvqkesHuQ6PxudLoeqlw3HBQfg8bzvU0qs81pZxcjWO3A8xFFhPEdt
pgHavI9KroyC/TnXOmxum/HZf4ynaZJa+FUbhKiev+G12Ap7ZA7ZnPgzCHoDcDLg2IoFS/QudPoY
M8WCP5tWwAGLOIUDxMPqHGCTnNjZ9+qGmhlBe5XIEk8lgYe8qHdCFuchYSeU4njcWxzHe6p8MqAv
yJbNYNy2AyiVPen+3enf8Sk99DthuA9tYPirV/THF0N9k+rdjjTrz71HvMez98m1q7fD/61wIP2v
nVbJ2syv5lsTNj8swN8H5zS+CC6RJ1+l51lg+Ty70CkCPXoXpz7mn4s0D5KK1e+AoruHEZlafJ82
KEj1ccHBoslVXoGkvd2vblGx0Rxmie3jhY4AcQWjPUpohP3qfO8ad3OI7ARgDvJA62pTrGsS28vH
CqkBTy9My5qeQtXZSCStcSyXX8gO+c77XVEUgNKAhgZuRbKkt9zJBdoQlKcw5AmjB/HfWhWZdozN
XGF5xr99pyl/S7fMQDLMWBvMg2mfMFj5DP9P3H10yXXuECl9MxA9wuduWkzvEXIwxqKBEWmWZkTR
OAOQefNk94xX5xk6DreJugGTin8NfdztBD13akeFAbsTwi4/udxxLawYjUDbEs2Wqr7JYFEu72MP
l8hZLMoDUCD3myxJCybRrmuwMDnIF8YAWvQ2nXoR6D3UkC1Uk1RhSEQQb756YkoddRg8E8oKe+2S
97JhNWngo26OuCGUCRO1QsHEUPnzdQNRKWuU5VyISwyG/OU76hPFiGpioiNIeUVEyJewNMI3MdKh
j5lVfi30NfUi21eGYfjPw2lsFYR+IlcfJr5bG0WX04jqojte15pNwQ9HAVU2NvQ5eUgYhMmvQi2l
gK1kvj20vNVdERymJtq6r429rH+zcua2SjIlMeAblm8aQ/TT6apYcp5I97oOZHaCVZ+KEWeCchwS
NOsRSynwrFgPxp058rVQrG1ho0t5BuCX8n4uE1LlLTEyy9Hfy7Yj/PsyR0gZhTNvQ+1e+WXxnpLe
+S5PBIe2lRGii+GcQYfxVolUBvxOlNFRHVa7/ver/y9UJnAjH5Frixsm8OdC6V+vy8ay5I5FHCBx
mI/6qCDp1PjN6FrqwzxBUQt9mUZMfnye7ue0Cql00EXQV3t9j2DEWuyhpqMWuvR9tsLicSIY2ZxM
ndO7CmJnqlPnBXgJD1OFv8D7BvuBNAOSwFNu9LpIghunB7KbetFngDtKPFCo1inMNIe+DrJqtSm2
JkPiRA7VRL5n6IwEgPLozc4RkTpXogOnybh8f2fiVCha3+cW3Ut+pIcLvKso+oTVtgsD36D2smnb
0yZ4PPITvMcNNz3NMNq6TLHkFFggEMnxaA+NKdN8l227plrobexqlIBYv+e2xxn3jBZ0iT/UwauI
YRulcCbZfwdzbiYjowcBRJqMg5NTAMaO0ZdngS2EIo8zXe/5yJqnAXhqhNUpcV6z0ZzrhZ+gFJln
hVjTs4YyeyadLOB4jH5uV/iIUmEaERD3hRE8pMRrPPLpdc+QmkX+c9m2g5TOgVHRnVcs+FTm7f5k
HPm4xoo0jCGonZtQVepSt6GmU3rbqxbYDxFpIw/RBHS8paekujgzNUKQ1F1FyFyznbiVCssXCObp
2RmwVSdM+ZDGLklxogUPLx9yj6oHNLblzEuEL4SszvGR8PVcvufXKwenjADEaQ0Nohi/O1nW71Au
cygomhKt+oSLroo8Pk3D9hPoqkjElABh+HyJ5KDsZGqdb3DZ2MWhOKvJjz877N0+vKnho/z/mXCG
nlZvSMI/5kCtmkx2K2h9at5k3Bs/j3NMcT2wjVunLH475DhtbqL0iT0Ag4TB1iInJ0Qv5E5ruo+A
/DXuSzltXlkbTu35WLDWqYGRU+mz5r13BJi6+bWYZ9j1qjm+OgDcpLDSBZvLmnn9tq7xSk4xUccH
acZipQ/HsIRpgrIK6t3/QZfijRyBXPv378hXnKy6TcQOps565WX1PO3kqzvzEGDwhPKWfW2BaZnX
ESFjbd0NAs26A9a4zoMjjhREMxhAbd/KH6aj7Mq6haK2qz/PCJidBVzqXCdqYkX/pXbURqSFr9eJ
aDxIocs8TNg0l/Va6Ba/NxvYdG6E7TC/75BQVD+QUCsnkokHXvNwDf5Rv/rlhLSEwBdXU8FngrEz
smKycMDl3jTAsmAdbgylgqRiAAi2a2ju0zv0I+sWcAFaz9EHBn2TRQEVOuD5MImp2CfnRWQ9C23Z
CyRXApX5KS6OtXKHhWVjNm7EVgeec52WjKy1yvxO50al1cbRVePW/ab1Owaasp2jxAmUQp0t/2yS
cwImh1tnbTOEhvp8KgIJjp2fk1TFvyvMdTjPdOdRTk/oZXGJFXnzqLQvVf5TosKxO0cDaBgZxzhX
bWL85s2Ta7jtLsLKL6clHiDmfR9m3d2lZRR9gXBAeF4w5vrUjSTN/prKIZcMjDcY91CcDY3BZKiQ
gNyzwXudZ3+GVgFTbE38WwH1vh6eHAoT+CUuvLKs/jguijFuxjUBeyKESNIg1YLhkBb0Z8vbX5Rv
i0shrJxF/uyo4BbdOKaGvL7eyfAKxbERz3NF/0TWZUB6oVdlDGwAStKMxbJwr64OEqxMLx7g8GQl
X+GUtr6DCDasuM5xCjAZGTsV+oP0FpXfUEvKyZq7Q4FRQP/ewkSf86fuyqUItGb3UGvPNHt2iZb9
VgJekS29YltdG26q0QKlPxnGZm3pU9acpAIrH/SM9k+wljNDz4xBprSXsnu/fBOsTYGq9lgW8Asc
Pb4O8LgDpmlRQJOSkU7/PPSl0bPhDeG2LjG/cr0NpzjCgvXY9Ou0ofV+Hm8/M25tajOD5SOXRPvV
+YA3cSzZy9EZRs1xcSpSequxaFYOH1tS99+mEbwEuHs5KnQ5UTuSqAUpPo1Wq9LgmVWtQduzwpwi
aCabpUZfw2nH3Bi015vhesgQTbRXMWazvtGhUqw3fFRYm//LXEAml0FhMCQtXORS7PZMvS3pW11U
q5FqVNJImjHn4+R2KuJB/28snG3g/FKhEyNz+wtL6csaRECRp4IvGFkyAkG5lQTF2SpQrtvbowAX
i4em2MguYpCiMHJLJp3qeam2v4bk+zFmgZ9M286wm+gKqdNfqh2MNxrU2Zozy8p1o/msG/EHYr0j
wTiwfPdE1dj+XT9aJ2Uhcf+11bnawO/3oLXaCyeVHzGD7T0TJsY5k4io4crvZ4HeBPp4BpvoNoY+
UmpWreHTvLp5J2uo7rHF0bRsB3OfX1fuqR0rbwdrAvwFRjV3jWD2QycgWLaHE2HRQDxxmsFr4Hcq
WlqEguJGS0s1dIrYW27fdJzrujcQTDCFR2QhLAYQ5mEpGElHL1OpalJ7E9sjjgQ9sFUwZVZH+s4u
3nOu/M8gh4JfIIXAEWh6uGdleBVY04Hx8reOBYubdhq391w3AbuwOpWQioAjsdsnaRNeOY5sOPxv
1PnU4UIz/CUfjgA1Nbm0f5hClGcjyJFxvTmRBGVIctCNZNshwwLFkfzRJFErINLM/QiAVHCTNiCg
1k4JXZJIFoe3zpAG/im15ulf3IVbtEll/eKw39LKfBILZx7/QBlZgXoZMFYuAzIgi4GYd8fj/238
2vB8mhzglzcZZO0yqWxplorbm4lP11BIGtB5SdcDHV1fjZwOLx503fZydFLzRxbQ3eYkTfhoGsQo
jOirDDmXhH6gu+T0JBwFwu0IEtl+8BRc88A5AjH58HL9z8IGAlmGB0jTw4mI2+6WlGmPK76q9JOx
eNTv3YItdKd/7wxDU1ca+h403dPaQWXS4I4RMW2iX/8473nifYKCh/USes2n+an4w+mz/K19nJed
chsZvWoj43IYS5RyZ8L3t9ghNHpP/SRrI/N5FHck7I1ph+sIiw254wLVASVHd/hwRCkIu/clAzNP
LozKj0SUvaD9tMW0BybV2H54cCnpN8rbIvO7Fa5PNs3UlMbTU92Op9708WZecwApv2MQHbX7DDMl
VtYSPliZP7ceo4X8NOAwoLzas/pKe/u3BYQmVaBO7O2YspHN3UbcEM/o0kE3CMdgFamGZVIKLdhS
TrfFyeOaFIQNnzLv6gij1yGecuj2Le64cgDpXcL0dftb/3WTiR7fNZCSKTfCcdB2OJxnKqI+YPLp
J2tocgyNIg/8SOOXaIGmxENGJ+jk8qkUfvpSIZNjt79QSRSGclCGHQPtIoMaKVVjVf+8D0eRLipY
xdvCu1NcErCoXUA6O7Qn3ryktbuaaEFmn6pZbme/vtc4bKlmo55c9m/ckBI307SxNggrl1Nns/Bj
kYZBDKbV+7aKqu4v083eZaszkDPMMFNJNw2beFQReCSZsEkpjbForIHjJolEJALbUAMrNLnPdy/5
dmaSUnGNtwosgoT0MzI4GPtwVdux/WkaQUQp4Wj9tcBAG/Bt/IaU3oT9puGx5vEHZYF6dMXzECcT
c74X2aj+nyqsrRXMNfww/cukHGK0F1w6uEvmOxTOf2u11fEYN91hFw3kNRwVarpNj62FuTyNbsfI
Jbk4cBGU+VV/2W9lVbrJ31KZoawzVkoXXv8NmdwJ8CQc5zt9KrlN5qvAeorFHqIPzU4GmFnMBA0T
nlA2xn4Wq6q3PjjAYmzl3QIfEjsCeU/uB6ptOZyDfjmRUZJOtabmHX3kNsXnzra/pfaCLc1TJt58
3MGrcWQJpqvc7T2MudAaFjausqAQhXeGAN04rs6nssucfb7CRlCDNghFyZu0ZnAp+hassVoKILpI
9vDqdFGMHm3mgzbRStyoW4gtfTs8I5fl3lZEagoyIogBmqJyNLiVtAiQWI0YhZ03/Q9xZpFAaOtv
47GitRNieLfdt3OTVIr/o/LTbrffqC8ggbg9H80Men5wCeiaENSHQ+q3JBCGSs3ZWwxtOo655C3p
CZxmEg05MpdKVvo7nAZgWbwDtXjGT0mE7nqlQjcwXQrhVkPFt05Awixau+QBiZTzUSLiXGVdvWMG
bOLVGnMY20t3KJprb/YzyBZHke5befcZeAJiZDoYE6qdYk1QVAjOFFCJdGs/a64JmEMHrLVry8FZ
P3D3kCKBlqZRZYC2McV4DiLwA+2EwDGx5azH2nlNrLsOUmUMlpHSBhtuYqkcBJ6m1pdVFkiXuXtq
G25R38rz4DSkKuczVXZn3i2i2h3xb8kdouxWB0zmH9Uh7PDY5venmzbxIdzSyKcwSwVZh7pQiMF5
guCgAyItifif3PBrMLgH0/4aavfpeunkMsmdXyekmM2qAKbZv9G8nPTrLzYWQUtjxqI3Gwwe86cM
In0oUuN1CY3jiZ3gLY835VJqx/gmPIXSODhRuZSvykmIOehClaBSPutgqcj1a4JG6NI8LeF7JM3j
aGc5ykoltmaMdNjUSxfwm/KebDCjk2S9Z6BRtaMZ3xdiPfI1OtlvAVNTrGLFJquRfRgUpZO2rKb9
2Bwzy+e5a0r2kHL6WZ6FAk9SgGfxEoCF6bjnzlNpPdt+ThbQEGULb5qJefqqpDfN5pNdxVUoNiUV
lAmUfYWHD32E0HcinWTmGeK+Z9U3qugSPL2nSg3x0dYuEuQMfS7WMFFfmQBIJFqxLAUR2H3SfLB+
gaoPW9dEF5xX9Tuaiy6iz4rHweiWnweAJXCmdypUaLJYKq02oOP0xYEdMPNwJlMaQVF7gyYX3mAk
vdV5bPEJyh9h1W4U8MuDL5MbQNIWVXKabOydR4SoZRZR0QU7/l5gDaCGWraYSJXjdzFAgjgt80Zh
eWcAxPJnVaZyoz2iRUeHXabTq5GvN9SfdOwM2bInAF90xT5w5hUlIY3T4vZnW544DZXI5Fm1yi32
p/PfGu4RABiLlUcQC7ZDLislyO5Zlc/Dx6TZYwTmz5G/MpbTExbXNVx6/stJwMejEps5GnlLiFKw
5voKDFDAK+MmakiDHTZOhzknm+XdodY4Q95d8DfSdXgRg+Wez6AW/ojlg8t9380AM+NvJZG164x/
/cPfe+xFdeBCz6LjmnETxiQgP8mM2ZdAZyU6F4D8Bz7X9qOnSSLL/23VCWkM6YmiC2EE8o3kw3vx
9uheApd0/Y8SlqZe6xTH6Q3CWAmv7SdMyE7A/fCA50GVjonvbI1bJ6Ked95SUtBfx3utVzNMX2Mp
mtl/8uH2l9/H2dhzRFOfLTl6Vc/A3lkU5ir2RSeEX9s0kZTAlPW8xUMSVhuKlGrYMr0bBqMjE/iU
BnH1C4YTj12gj9v0+GxbsYxg3oJlUoQ57I2U0NGSsKh62XGDa9cEdCdSAT2neIkbaS6BGkucqx+2
j6OvvGuO8JGUvs5VTWFQRTp378Q4PNU8ELCNOE2hFDlzaoS76SdV1OiSsunbRZEFU16jrau1N2Et
IcPAGFDS6T0Z+b5/j/CGewK7v6q20KXxmdhhz2pYsXkizdPtGbZ1E3PxDEhkWYzv0kQbDuNzkbkC
FOxs1nHeSTn43cPrv3CmPsFd0rj+JU5OqXaBw0wmedgrRVIlO0sxobfUtpcM1FDu7NaGzGrB3uRF
a6WgHg0ICOhA3L9Vyrs1TrELSPA9lni/L5wr9GzOYWI3ve4w8sqRSNmockpM4VfaA+rUAo9Y9OLZ
/JJzOFY8sk5yYIcVE78q9NKXoZU/gSbrF4s6L+rSIUGflQjWOveyfc5feaEFg2U0AJRHsS3kKzH/
85IdEjm+YTJcslTiGlr5Q/clb8Q9bSdkHi3GdprulNVT3zU3wEdYPY6e/hvNVVdGMY+kAr2xAWOa
1yYuMwP5bkK0gYSeRefU8Cl/wRYc8bZdL0xPRuKv7Z+1GiU4u6gbPm/weNSIJhN7FkM4VSFIdrCN
nr4VtCEp/3KMo6qrJjKpMLIpPWSdH4psbzUPHfp3baTBzzVl9JE7VNSNMve09H76Gg8MUo8fsKPw
028hTZqHbco3UZK87LG360SgM6yGtD9jIFJguvlaMFhPd/jExnDyorxDuRuad2p0SrfUNySEF/T+
skft9ALgeqbsEudI2hHRf1hjpUf3p4WZ4jlavyuwZNV7ABV/yiljLvLCn8An0faPiYuDXbNU5cd+
knmjmG/D7enMkC8OCrlTWGsiwgupuJHNkn/MA2tB/DvVdOpop/cRWaaABwvF7ZGpNNs0Sb1Xbiwr
dhz7sPTEFKSz2+VIMIebL9ycOCa79kKzvrzTiJUMp6l7FD3WCe4k4WBZ7+uri63tx8tOUrs8FevE
gjpmhmk9V/hDhGi6E5dgO8WOhSgBIFU3QA5LdOgxabym8iPFoG8F7f0XG4yKiXMwOjZhmqsIb45l
xlIyJZDF5JBf2VKxt2rAB05mUrRTPx0rX/eREzwu0LDSzHbua+MKUaM55/sbFgSORaRErb0fIlCm
7771wws8ut0YzJmgH1+sJRi+/9gfCRop38T9VOD2JZNldSdTe3GRZz/qgX2OVIy/QneJpRE9Ctea
ZKE0P7ceRA3d4bvpMjOpC5WlAnvXrjNSrZRNj6LjziSq94TGqLMLMeLoSBPLRX8/V4PxM6/uQWHi
U9S5oXjkGgkR8SDzHDkn1yuyRwsdhE1FBIKPCsHfoMPqOa8Bl7sjGJFY/AJCTlF/c2N3d5G4b/yZ
LCwdYWuIg4H2FstG6CXLc6duwxDBB7inTeZf2H9OVubJDvhMSm3a0wF298yfzVq268E41lrU3vkr
EA04J+/UBv2n6Ld8XMbLqFGZ/1vqhqzZntLkfhhJ/MuRR+p9Wcc2jMWO4POg/FpyPhsm4QBnvLud
3CkvRmgbtBlE5KkWciA41xm+GOdWA3LbaJVR+UtCsVQK099/F3QwQ034GqCTpB69+c/dztzZNMU3
8I1YlFiG1APEoM0Wi15z/yr3/oxG5PD1ivE3TxCoFhdg98/EQUx0lFHrOvJ1kUK57Lh3W64L/X6A
ZWLtQiKryU99QCwkOCbNVc81LSURgJfeQO5rOR91rXYsDbSOOAl7UtzJrtl9+rKgZQ76wGhlFtuo
mL8lcz9dxZYI3VuHzVWWBc7mhfSAbVXReyWjmnrOdoPbPAL+PxTQiXmQwfYThLRGfCNhezB0Mt17
CsI+oMb88LP6R2HlMm2OfhgBrnQA7cdNSDolo1dJ8/oSYPtR4GfB/WWXirveXJm0N0nNKJamgybD
CugBHEVcgKgq+thmDiVQ5+wiEKmri1foaviTrRQUh8krAQ/uNCkq6EWzoUBggdT745aslEtESoSc
o5jeQUTo8YjeaQ3x8WR58Vh3rkzSDg/TDGbcVYNvS37FsHLyY+uhZ95JVD0MmDVE3J+t8Cej/v/Q
/PoHvUyk+0W26S2D0dNEMMvK5qvKV5CFQUL9Wl2AhrILq2uB8k2aYGxJeuz8u5ylGLN8n3Vrg6c9
qPV7FGytuBrBWjH5wRYTkC7bPn7LP1uIEHRZUG4eLF/ew2SXk3gJprLaPDqQllzZRPoIVwVQJgSr
QQQpQXy9JuxzNHXZFQaBGR/9iSFA0VZkENE74BopBjs0xWE0k1utX5D43Lbmr1kH8biAC96uVE9p
3qIUmcoS9J7Fcga69c4KTdvMtFE89oWWH53yX9Deba+dJNDPdHOTOTjYORBTcpZfGUqnmvU5VCo/
VKmovW3On2ENqOdsHSAryrboq06vIbqelqQJ+sDunpPd1EW5NKTQQqEJii0PTF8soLDZzMuUAvMl
23OtjqJOn2H/ZVEcBLPGb61TKtYVVb9vO/bi25QqRjzaxwGds8wo1dGD5wq0MoI1EL9cYoxVlnos
4JGa9SAfVev/Bk9qzLLbAB7lLdQgRkZvIabcd8ScsUKTF2XBX/W9b+HH3c/OBP8F0dLnAb+MqTJl
6Ea+857dFmUt1AVOuPqNCS+j+GnuXPnFm3Nec2nmCzohTtMppob2cndVoMpUMyIs3QVA2hiPu0dr
hC+eVor62qzvZSjUgf+GhokNNryaeKMK6Tl9QdypfGcdu5+qXohGNz7GAzuEiQFbqeC5X+xO38W3
DFwqlCv5RUZXjfse2uQOKK16XFm6v0xcznEldjJp7hN4WuzBwskILWjsAkD7sBvNKBQA/OHLHRdU
SdVPTdLKriGfU7+gNg8Dfr3PDLmd3pwpPkTHHLaribiWv7nGldj7402LBKpnLwIaJgeqig7pXH3a
2Om3scZiwc5GBoPxQxoDYvxxf9otfg4FclXW80z//+g8dCYYQqkHM8TeuMdfp/IBBYRQvOXWbuug
Gy7OS99UcNbXemGcCwdOisXufuyyH38bo7h30IqI1m/9GVJlMI7JkwpVyfppd4/Naivjxvy6/K0h
WqfKqp6hoeYP++HaqCLRbA2UdgZNTs2vhrc88RmzTIwCRWScbkP2O7hjtzhXrMN1BNz04jvzFMnX
qoP2W3/NcIpUzk0I1MK17FM/qOnSG0PPh0bavzH1roRz97fpHe+ub3SRQM1E2N8lz3275QIMFHsP
r9VBW7yox97IGviOVzFiOm2eKomldtMziMBHo/+DQBUaRMT2+SRiii92MzIH7wZ9s+oZCb4yMSHt
+5kLsNp54wMnahxcCHyOjfVcNlOUSH0eXxWPofRMV+Aj6z4RVjPU2B3lYi9I9wsBFSZhS764hpDc
drhca6bYsw339zhXXTMEiQTZKlmMm1lQ66luTq1CUQrmuu61Py1/khrYNA3LSkUXgmceTSvHOjQR
bhXjDI0mTWstM0V2B8eFlu5jMCqn/QeAU2fN94IMpq3BXz/2Wl8zHYHgJA/ms4MqPWaOjM9ZG2eM
gOs7K7O1uAqtKnu2BFjQ1y3qzX6kBe7idijiFuotlomTEk7AmhOIykHuG1nF3F9NQRrk/H3vbE8H
Kv24WgoP2We5j/WvZSj2j3uvsbWyxYa1OliItsp/6UwnchylXfH9WP9HNnbVl3XbqDHJVZLcze2i
uyJbpV7EudtLQA6nffCCc/1aNRr20AnzF5heLq02FJ13HqviYbqHuRgQNCMSj7zLM2z794mjvW/w
dzGp65NHM+4LK3xqtLPg9AZ1aaX6S32yPpQ7g3dJ8tvtw2RcUVyQDdQU/x7AmtHYLco/gIKU9U6o
2m/YpDx0ZOXNEOS0C+u83Y1P0WtORQ4TKQmS+ZGHT9jhZp3Qb5YSDe+bLLQKsuQCDzW7DnsxiAN5
xNsLAsyUDz8jgt2RKE1aP7Ad9DN+pCodAbCtKNaNG1Nw0h246LxRWZRHYwb57gzeJydA4bsRFyNV
evPh23mLKQgMvpGQTZQGKpo7jvlLkHV7PPYD/awuLr3JlfKQHok4gbn09b671kk7fXkkS4Td2b6D
z1yRYv+yzedEhclBDy1bVqTpnAo/T0h/r/bBNZRQzqGoum90+sCSdBq7Rsld/PJvpifmRc8AF1RG
X5v54GoTrLhLXtdvmwhgjJx9mjVWfMBHGDXfPEhMtBk0qYCWwKfDBKyYNCOnO5k8ySJH8+xV3gIn
qzbH62IyDOUQbB899BvdtqSph021d8duDlZKJ7l2HTTO6q++QKoQpKIZ/Xy0UWot2CttzoQ+2j53
FsxHxx7SsVa6MgkN0FY1mgj5Ry1XK8XGpAuwDgSg426U+VyAiezESDuDzvta4/Yt3jTIKESOtPjd
bExDYxn244Q9W70FT5p1Na5imP3pjjnPI9rD7+3ldWkFPlSxLyhx+21uJWdp4i27UL/HcDNGwipK
e93NjfF8/5qWDICbvEQ/MPHwA0otemXzraj3o32H/0kFBKMVu+A0x9SRJMc74XNWSw934VbFw/zd
RAwttO1priziIohdkGU9Dq1X2mcuHa/NQnnKOiM79eyxwCeUgqLk0Z+OkawuRbD0kyoOc/y6u3P/
s4R6rUdrJqKIwnMN04EnWnaWDtDjtZJdYbhE8vspZ4LJ3ymk/QNDejFytDSQT2Dj9Gapzxe+IgEm
5bFPtIv+rZWYgeyooqIbnjIpn3dXkTvIVMQCC4zOO851XAENciu719TAhIsTTw6DTRU81JEiLAxj
SiDco3kIw4DdJREqEkajHp2VuSCG4YJRjf9LivyvQYcfqjgwHtLLOuWFyFxvCprFfU87krhH0YKo
ONkB2KLed00LmKy5oQarTfKk+dHh52eydM6UG0Q3wwUMRgSJJ7/b1rK10wz6TXWHyb6JwllE3pRB
s0nsn5JsGqYVOdc9aiF0Sklhd0BBOXCYxzqqLFeuTxg+uC/g4CR/NCCSPbxsr8pEJQUPq8AQH/8m
o8F3VpJW+3R5o299XQ8RuiunQV/8FXu0GPO2hWHU15wPcH/Xa46YFdodRpzcxuYt8+6a/ftwxLgN
cwO+amyO9Bj9LrqgcoQZQuL3PsbJnQDUYsbVZVJHm3g716Yo05bbssP46Va+rPExpuatBxUUjVGh
7OYuDWPo3yGEwF/QAqELNjliu0ZCdERhQbu7hKgebXI8xjowjaNG7JUmdRk3KwYlcjl3Vl5MMMIS
NPSf08sK37/uC+T5c3mAfXXkwYyEoS4+ADYKBgp4/wWR/CSRF8Z+SrpFRPS2MDgYYDahxHfFUkTt
3BlVhtHbamcr0mvTSZtIOvgMi0OoJPPEdt6h2/WwKhpShBRyU3Aq5XoPh2Tpl1wH+v9rxqiDl+vS
qjkv/fT4nMQl7s+F9L8QNuBgWQJl7gxHaFUuUvlHc9mDMYSZTZQjMAT/3JoNw6JZiAom4OL6/ayt
OMphIQKpqNV1Ehnm4pOvkvfgMtlNaAz0qVtAeuypsoTnzXU8RmYHHl7i8HsWM4wHGGKy4MwvXwJ6
zQvTS//5q32UPgsRrdBFuJNfW4uFS44Sjd+ahgpmVguKilsHXfLpewe4ZeOUkz86Xb/Kp5P/KDEQ
vretc/bSVZfnhYYq8Up/hEFL03zJ932CqFmtc7TYKE+b8ZQvmnQ9+S+qswTTF9pG55vmNiBEgZoz
SO3HKaXQBxzLxCBucVdg99Cj4Akw4mNnz/2dcUPG2UeayypcAN0jFMQL16dFLuMVfxAStWSIIVr+
t32ugW0ZsrQjxjqPUgB7MJlDzQhMlSwSY6T14B6mFy93ea64kcATLVtSlA+GUIPDTRWfKl5O/x84
Gw6+fd4vcs9e6CYg+hnIIE6Cq+/X3Luu0DFN5gzyPLAGpukkJk7Qo7/rgnXSmSG8eh0pmcWON5Ob
blj7b9xSIvexWA21rZRDTEPdt4A0PKWOQBEswwuZrVhdOpOXz0aQxuMufUS7xL+6f9eZMsi4M9E2
eNFeF/VL7BjRGHO6HGtVq53fbqaDmfwc57V3zfq2WiY8oUTUalgCZ/kryrynQKJ/D6fIQuG8lsAD
VQ8ANI8xjavvrnSZNSjPVrSvmwWszMpYp0O+/hx3ORXMLIQBOhrc6s8g+1VQqORSq3thJh4JHQFm
MRQYMvAxUbjfwAqGJESZ+QtZ+M36cVcGA++5uGli3fwgNjYTfoyhtc6k0UFyzmcawet0PgpsB2U3
mhxg+L6wpCoqyF6h5NaRzpQO5afCEDFV7tfUZnVm16htNQPjmf1sj44AAVVAF8ZIOyk3jG4zoo5R
hry3LrOfqP5SS0t/aJxE4/t1ihTQpV5+YVD0S+dtSPLyIQVkn5EH14TwXZc58gPR6Z2qP9vyfl1Z
d7bvSM7O1bonGFHcIZI8txGmz3eTYj+X2owF1EReYVD8xQOyNatxIMa+VDgYiA8Bh7ExvODm3y9g
Qr38i4oMrved9niOPJVTG+cW8EZRYZ3IYYxkTEHd+NasIxgeXPhs+L4PEk3BhzjcB781e7vNPOxz
DMUvKLwhbJV1pmRmETIXtv+nXnNdsu8JCt/DhPt3wPQ+rQUyuhxJq8Y+ykM/RAvCEuk0jw94IQQN
ZNS4YYoLQ+zCbZM5mLGHpH0mrwvg1n316c+SjkOxhbGb2RQ3ovsgSxW4X6anBwwINiTYAWrfkTJW
HhBfoU+PB8Stb4SKVIx2dskemqS+a1NsbKphVt196pRpdMSCT2T3sw8RHFwJMs+Pj8/oEB4DtQmz
VyF4pRQKasJF2HNadXEOaOLw97neeexjMP6VtDJdNkCrXIC0dAntHe4zpKDeGqFKhM2pVpCSxGHZ
JKnJZdZkw0SHLUEi+xAAJsaBZaxqizUOGWu/DPBmKWBDyZWLpj21l31ruiN/raP+KJ+FgajdLjvg
unjwCMrs+aKJVH2PyMfxD/ym7/HP+pvJew2HWg9jPQOhPyeKRkyvwmqwkjOsEHGQLg6GLqI3OdFz
M2tott4l5eVS6PZa5sHpyx+Db18VfvjRecCrycTSCUazB6+TV+9zv/rv6kZNK9U39PmS2F/4DHLH
rcjA03iAN9mrHJ+uiwrUuO4sqxcIhDk/ro3WZNhB7gVRexbt2jUPZPQlqd7ms2nHucDzYG/3Kb0l
M9lVCK4PHY16EIAr1MqA9i4q8bujirkIYYU9vz/YAfgelt/pml17a5RiXFtmwdBkZsCSnTbofdqk
XvJZU68DG2SWC+wY1w8r5SLDoYO1P3etD69Q+ATRWNv1vl5pNgVynI0sNkUfM1r90S9PU+PhbmWF
jz33E2ZIyM+cuH8m98FLe+l7/QwA6pkv+G4UDfe4oIFbaL6yxTI9P0mWxMnodcShg6cV5rtBPypq
6yrJgyFBJ/8gv9HrTKYNSyadf2FInQgK8jPcE/djC++4VXC0wpDn/N/SQUOLDrDXx7noAJkvVnKG
XGdOrwVatJY3IrH/6j1s3MRF5eJPpid8X+J4Mr1DHhE2LB9uLsWCMv9JH3Q5eBwW+F25ybJUKSxx
ZKooSUGvaeOiSTm/37vc6buz38QHecY6ewvbpvywDVVcX+/5qXb3TdR7snNF/9f+S2GkCFrZghW5
hrstekRzNvk3qUgaLaGlGGSh3HLt/eAWYpfUYniR4RMvgoR1BXxbHwlG//dw4Vegdm9Jcdlb/lZc
iotsJ8LKIEnfORxwgc9kJ6yhZzkOo17+G8uBnIqZkWfbvLpePqT/dmVpU8oIepNGfWKTo9xEfFbd
Dp83yOh5NhiIOgnar/E/Tx8e8CgGvEKY2lCZe4RR2cuC2HBQFhNFv9AFEVzY8UWAbsxPh/kbyoLC
lYplq8bjQfhv2pbNRdzKyArYeHm7pWYv1Tv6JEvPd+kjcmBoIG4XrNnJ3rcYO454UAQ8cYjNJjPg
X0UWuVZ2Jxm734HEk/yWL7yQ0WqmWvq7OKLBm8MroL/t2x5s0lsCSe7nT3/+9nf/Kcq2sMRPjCMA
JvlETCgjJb1h3aFE+dJj+SYbe2pN/2qH9OVjY6gOsKtceiYxHxTkkbQJFXY2/QqyMS1Px8iRUwZ0
eYCp7yvL/JgUbt/NTKmoxKejMkDNsALpjnUu4XvCUK3pEpMy7AUQ32xNwxN4NZ8L/WUhH+XGwoba
dAj7fJau2otak1RvEJh7x+5r5lB7G9flVBHQE1XhnGfp7oZtQBfanj/VldZWtSDDYe6fSNHkJMqC
QgMm1KxxVTcjeEnnnM6XFYw9pm6yMeza+xVLRSQ4/UhdRgHDeeBSymUXruX9GaDBSOowPFJCEGBD
6pVY9TixbskdktO/iEsPQmqj1RUCup1k5TOoavU22dpGTZ5aWeiOurckrxV3YuQiX/kwnc87LX/j
pSWxaXv+sL4f+iRG3CQBY0GeWrxbGmlAwFsHkUxS0V/9OkkuTj6y87+psXdXHaywWOvcYIDN8HCe
KwrbuaXzLks/uXptVaqDVkpXiCFeeEp4yGKVxo5wZoyJkkAuwhySoIoHXETJt3u8Tx0IsrQ2lOmu
zTqwBqs6tafxFHgDem6OV+Qc++pYVNnahCp87DkWmo08TE6ZCCxWfPidYPGHZjmLqClnqhbH+uT6
AImtpCYhZ/NDj0L6GwPz/WCRLsXfPvaaPvLDAgZHL3CF7AftYrcjUpnWEH9AJXCA7UFR3B+4l6Ny
NBf3RZRtXPjXqGoXU9NqA/SwjGT/z6bekmcrZx8s4ovaeP44cYvRdWMp1Y9kz7MprmzlMtzwtRcD
T003hRAxIvcOOsFQUhFKUa5Kh36zHvLMz8PaBdmN+nI+x9G9SAsz6uhwZNk3TY7dYV6UP/Jwegzy
cRSxAcFJCufNNIU9W3AxtjsKiqOrk4S5O2NAswkxV5D4dwxcDYcyjYvCzDNLT6XtoX/LuGgwrozJ
OoeL1P3xGC5tjNZDdRoehIMjqFWLenGXla868YYgb9rMM7BOYJJAL/Cxy0ncu10AFLT7U2K6QkbW
O0MC4pa8qFNu99aWcAne3OwVNChx2eYFf1TUgoBcro10mjpnMpi/L6GxDbl6ofrannVMqTMOJjCN
H/id97oNVGeFNGLuYDBPmqTq4BCudgjd34HXII+h18CjVikZ6caGJKt2oUeUyyNpgBiuIi9GQfRS
Npb7LGRuQTAG2khlgFHdNf1GeEczNpz42lnKNhzr2zLI8EKW97RxxnKyLmx9dGbHR7McpLXxKFr4
UC4jpekFVeJYZ5SK4gbh3zmy3/uI7fZnerz+n9QBu+FaTHWfWZFKzS9ZXH75zjM4KIft+lejKxL2
qP7FDBp0WF9GSBlEpsVVZ1MMZf++8s/mTCnu8mSdU1oOeL94TAAgWTIEPEkj3ZQ18yoALhGgtbqN
27pw7EWPnLNTANZJmGKHCGtyDnM0bEePrZ5DuC+7xtLOWAWU9e2uf7nP9LTdRbK4fUVqpezHxh9F
vRvcgGMS84GURLAdpXDMQM2G/uaTMqGOmM+Sw1wWxNMB0lWvJ9d/s7YYVnUz3CjThG40bytSskSY
msJbREjsWEPV7frqqZqEJRutqIO+U955G171CSHZCcsJlymo8Vkuwr7vNtyeuUNG24B2PfHGlMxs
AUIsLSBQZY09JIWAmVCj5X89Y5vrjDMpBoLHNWNaQWBr8kTLaGGHkMlueKGmXEt5k8ARt2kbELj2
N+KvLI+04/MkFtdMWLmHQfm2Znx76RgZOzybcYmonrBDML/d6yR9O4CmkwR7CUepoM+L6nrOVKE9
pFqQXCI0O2JCbdBMmyfmdLsBoJyabNIAVCIyzm9y54uO4nUXgDHkveIzG/IUqxYbDSFdennZ3vTX
k65Mr01/P7nJ218cTOM7ax0Ln7MRD492eWAmwBfL68PnBiWMLCqaDp6Ty1A9igEW1gPNQ/fn/IIR
Ac5/eUIEL4ZgnWTrgzaE79NoI6hOH9mkuVdRUnWfIdATv6m0xkfJl4j1WL3eIO94jlgd3k4yFtgF
v1OvKRsf0hiBMcrNbollGZUt7ucfT6xBk8GL8nulS2r8Z12GRZ7IGFsJxWH10K/U5imjIAjSaNRz
vh5ssLAKbvLhiDnZOtQctfSBS35l8zb/zDAVb+NNFNuwy8Shv9pIgjdJ23UqJLyKKISycMTTjBzd
wFk07efDuxmzwrqAyofkWdg3DKPXhjqUtEgi2bFtAwtu2fu5eLlLXRPkBycb/WVTeR3bFZGIbH7W
JqCg5rlHl93uC58kbWyW/yeo6B+0YIWP2lA6qKUqBELpN9Y5iQNFgbTA/oupeogWH1tSKjXPUmK7
mtrtabW+NzGB/1AqVktY2o5ympNE0X8KonSper6viKInZ1gD8F2JfdW9QTKNfe/8VlrHRn8WevWl
cfYLasynHR8+zqKCP9wVCAG3sdSXCoq1HE1XIo97yo7zHikvUaz6SmOhdMoTjjZzR8k1ZIwmpQK9
X9NETxkGU43W1wG9KcJ2z1b0Y7rkg4P7KSjPeV7UETHmgjhuz4UAOjuRXJP4ZKv6fv998tCeWFUq
kY9cnQgD+TTiTe6NObEV5iWK+CGLDyGjyulC3BB02aKfWvUgtH4GOXVYWEPAE/D0j178HG36hJx1
RJ/fM3UiBKr0VY4e3VH+puqqvlR8QBCkGl/7u6QcsL4dG+zzjAps9nTXNQknXfkPw1HNR8YALTRU
Agt9SNxZhtbaHOu5D88vA7KmWTWG7TSAItQrs0aCbxlGk2Yy6cDkOU3C3sQg0Z3oMOe9V79rweMR
8pyRSemXBlsv5C/nwDEoIh+jCw+ebanP+WGqYMGTm+BOWFE8bAMayCWcGmt8kG7JO6wgctepXBAr
gaOk2/8qvXSO0nyyE7mK1HTK1Z9B9qEp/XuSk1HVEA5MJhkTWrLt9bMzS5p+5//8TaKmbK7l9uTS
o7jPnLT+Yld77sge+2z8BpLiUiQVOKWY3QHjC13MPxE3CXNSJc14DV/4MTNJGHA67gZLbmgtQ2Ip
GPYRQ+dFVamXIQfGRqVxoR4f8dmca+PRkfFcufAH9r3fUmY1h6iDRjpPy1J51gJ+lutjgra31HoZ
RR5cQNRPnKNvGHJ3EVEYHloPD00GjqCUO45onoDIi+gXvAFGn/231n9kjjtip5huEIu9ZWPlqHu6
ytP5Q3CGU6Y3idHEEYEhle9IuYQ+xyjengVOHeg5uhZoS7B/OPD1PtClpE5q93jnbC18GoACuyVo
AlANaO/x7L3hcvJj3OzUkLrmK0WkQAKpkFLnXtqtsq4bHGBmIQZxI88/MM8AsDImXuvjuM86d/w+
gE4xHpixfd1DPzS9bSWBrH7o+RYruldUqx1VwPm4LVe9KS6AU+CS84cgoot753M2aXqwklEzYqcy
pC0CW5T6pnffr/kW54dJJA0oqz2x0CeeYf7sircX0W3rnb+Lcf0M8O59imo2+5eHegSaHxPNwbTl
/VKiKUOnyuVLmsuWQ5k1IRY5sXnNuNVCOChI9IKIzScZlqMezlOVQa5A1XX3lbo/tepsfrenCtiN
MLjGjgKwrCKhW40mlNappTkcm8H05mgqw34mdPSB3eAXHcycHS5DNjcpN2FWY/NXFyQuzEOtrQ2W
SKu9BoQpp3DklN1k9u6L3zMjLvj6bhFyXMS01knm51DM3ET9Fap5NQLhvHKSqJzbPnaVqkHECjjr
4vmmyPk+wNi3cVVA+7F1qOHLak+ZZ7Nw+MlGP/hK5CTox82rtGm3sY6rfYzPHmnee0dSCwwiiMAF
gaak3fKeGvoc2Sg70tThy2itY+Vl2Hk1Ocvg/MWhgFdgMESbna5C4NfeeZ4r8P/ggmhLluVBJIlM
pSEOgN9Jci1uJXbZXzkOcxSKWWaL1DGMsoAXHMtadKFXafhn+xZAb/5fGV6kTxYw25oXlnlSvVA+
Wzb8HcYMb6FAOiXa9JIK1dn1G+3SvvWscZ+7ZRD1WpGgjbkPRN139q+WDenyjZlbiRnd72WYz/Dt
1ALOq4DXt4QeC0Dh1s85lknWJT5ulXxnaOrDVYNNnIZ0NDj+tN9y8RNtUqdqdvG3+s1Gax+S70D0
WOsT7B3aFILYk80nbSRS+sWUZUtSZebeq0zvTCwOEMAcakRppWXXFWcb40YWjQzLXABHPiZJj8EC
Qgdk3xld/TUf6xGew2X+klBIV/CfaL7X00OiKw8b18k3vX78ydaoPgZjGDX1E0fM5G+raPALT5tW
CVjNP08+RgcfrqGKzm6MQr5GC/42ImCs2Oe1YPeV0ljV3iNbkiy7hAPmvCXmiy3sEUpxUXpF+v0H
y7YjBAEWDG/haQUqBvtiUfmSn6GOG+Oqq33oviDdKK57JGe/zURozHccfsGdjKyBCcSvIztOf18+
EwGoVuuMsjyPEW2T6VkqSYpQhIXdlX7dNYlQjIvhEb9zgWJOUn8j//tkqmFjcMQIgb8MqmoEW3+D
QEHrcBK0lDSnvdHxUvvaOF+Cz8MaQ7OnfSvtMaNzg+7BUfP29jcvj3ctOL7L4b4KObab7ET8pUeR
nk9bgidY0QAbisScs/d7D1VQEPI0/t+fjDm0bMDL7sjO0MzqC7geAsN3RNWLKFImMrO0KKvtMTZN
h8KFe75GkJiMIcY92XYDF86pNsmBQ+u2NJ4eQT3nlQxcpoxzTQguuNSTG5ZijWtqtrPFGMmQzaoQ
HM3XDL674cHmTRi/OTkdkvtkfA4p+Y/0fSrD3SXem9z7lkuE8/IVVAWoZ4gTgP6jJrjTA/69bXAq
WgrawsvimZI00ZvbCbSZ7Ak5oDGcQi5Z1MItqljQI+69s4zA5H2IGCLaMOeKMCFhqlB6y7OH5GbK
I/7/4qdigAKRqLqIawnyTLtH8X5tkDBH2ehpaH4/n8vv8vfMGRfcuMBNN5NSFYfHeZXZ1oVa6IqY
CaZsTJjTCPHaUwY96C/t/kH0b8SK6YqC413CT2Yj0Q/lmPl3LyCD6+PVZxtdf2XbFB5XB8pTqNrC
Uzfn+CQ4uzyFZVsBra4/K7lQ8zw4n0zQIegFdFpZgEK5VMjKNzq9m4Pu3BDUZ5nOs9hVaxGl5RP8
MzYOmYh4hlmdh2PtgoE42KLrTUAbmri6Th0fgDMXaKWDA3jlnO6ooUJl+XCpfz2U6a7bgn9OuS6q
++JkA1jI0g2yPZw9JQOuIeAEDARlx4z8RRyOuR6xlY8o84HiDloYm7cWnuak3pN6AVZb4GgNxrZ/
DxksvaDEzg4kCzcsV8IlXvd35lwKEfXD7X6Tt3Kf62nXpEjcHwRLRn08CLwdzgyUeXVxm4aqdYRM
4DWJH2MZeKXk5TVfAwm8mm89vfgItmmu6hpU7XPU7f9lVM+IUpCUQVxxFZyEPZ+rWT4zG5lmWOaX
ZPc2DCUEQU+G9DCxCq4DNQM03WmJaZDNZ6Q26tEXjjk8aE7MuWXzd7BV0/HD7XWJR5U3p2XcWKKX
cWQTDlQT5tAndmRRDd/nNiX7UQOmAD2zZ0uoJxrfxDmSX6wodZJJc1H2i1zwmQN/0GbxHmQFmvkq
4OG0kbh1ZwHNh6nX8arx6x9v33I3jqRyQIquaWgexft4TVLvT1cr7pgMiZRdtg+IAXpVpoDaWDqy
5g6HzQVM+xKlCVnoqFqHymcQFi9vb8pGyef2cMkiYyuEFjzxTO9q8TSkbNmiUwiH1om84QSr/XLb
oW7kPlJqHlvB77+q4kZwigpP7qHy/f/HPq8Bg3uZ/l6Ft+bK66F8tBXCeutC65kgn/Fcxqwup7LX
EIm0k06S+4gkUYrDrdODfz80lFdMMuREZ5Y+bS4OYBALo5U6rdyjmZ4ng2LH0eY9ROo0PzzFRAfJ
v7VruGd45exbGmTqpzYZAik+s207LnavXswEXatKThORMQZFAZIyNl0TFrGGzSxXCQhj61drGi7h
A5ePjbhOCyqgRFwJsbHf/2Ye55iIgajPKJGB3IHZOClE8TM2dPTt4VvtxUGko9cAn9foYQJAkiVh
X57YItzfsgvDLA6vWXBTPmDXYCYRiG1KsUKtubuRpfSJgR2P0OU5Q2r53aaGRNhq8MgSM7lamft6
44EWy5O97hFf/dP6B0MSF1Ta2aFCG469W1/kQZ4GI5A4zgNaX/HxCMdtxauxJO28zMnZzZDxyja1
PASCdMB00Az9juzYYpm/KWhOjRuLtnO79n4FMWFQIVWT9GT5ZdV4OE0IjBV5aKVXtVjIOHmbWfeG
jevvgWRFKwk2Be5AYl2d4X/WYjznloZKws32UjcE4VDKChxUGzT6pjgQRZ+bXhHtLaeD/sM0VFaS
kOK2mEN+/HpsVik7irrkts1gAVOmzug2+Aqcx/s3sP0u/UmLK8XAZeHunp0dxaycFH+7Pj0GLQp8
BAoLJJIBLEJLMcLq26ZqiMx1gHhFdswm0ra5LqE9fE16KApFTb0WpYKkAE+4DYCkL3RVQ3mICwz/
GHJiWE2XBr27l1dEJRIH3h6bQ1r3uKcaPHRxIEvbEt6i2mmfc/tng+PggPpYLbF2FwZC9Gkxbn0L
I4FKmWXJmTxnYIRza8V6/6iwvkR/6+GfuzRS5aQ1zB7SGaqOzKn6VwxLFiV7WXONM1FMrQ5m/0T9
lRjsZQhP8nKFd5J55zqvFvAnOmSjOGW6QKk0ON9/U9dGeZXr/TNFNW3O9BFWtvt+dCr1XEHutQB2
XThsybQJUodw3xg3BBvh8GCLove69KnbOQgBxUzy03cvEPJurUT1LKMnUZJGvut+JGXRhKWCtrkg
kLiuIWJFjX0Jn6DRH3XXe5/Z8RPBdPMc3ARzddMuCBefzTQ3dpnFPGWA7fCkrWTFOkOVwdiW6VGk
Ty11HwOsUTa0AB/KNPtnM9cSG5IucMnAH8c1PiHCzsiGe7pwDgwbPor8hfVu3C4+rvwhnV6EMs4g
MdLiCCA/WIU0Zme3TfZ3HrWkn+hbtzNJTADL5lXWzGaSKK39LEG7DK95SbVmXOAl/s97HC+Oat08
VXKh6m9OYvwIWEirhYrtuLWLOrCA/CEPMNjVXHULFNnBfFUyNv2QYiATX6hQ/UAOGtT/l9ZP9vbS
KSHUM8hhQupMhWMCiAycY3CnNipX0JTbqJ1aW/KrCy/FuadoWO72QMb7t1uTvSrDGaFRWozYZXNQ
ev3UqZsNwZv4kjlIB80m+IWdSL1b2nzBoiV6suQm/LhhuF8juwK+NzRZKsbl5R4okWkdcRcUOCog
Hx9L+yn4QDKnaY+VAh7mISpdHh+UXxx33zRxoQV5izlJ53/lAl2ELsErfZY9DnJd0+Mu0aBBUMYq
cl7p7Ia6nkmrDlrSeMX7lIcBnMnEZkxeGez2Dc2hvZks+J3fkh+ixGt54fnvqceu6j6+GbZWyAeq
RagmrCrxfwEmptdrz2YsD6F0we4nvBPTecGvtHDJNh/hVHt51AhPaGOTc3u2ItoY8JRWnTZG42o4
rG84WrY7/LNfBUYsSrPzhh73pSMyKw92p62TwUFtnq3oy5IGOXT+3XrW4Uz+ZEJahJHv3pfgqBZF
Vjh6y2OoqXZfQle9PD8sYHbJOeJQYOfnzslmI+MaKdVWx7A4vc5tot4NFen8j4H5N2SMB+6mc4Ri
3Wg6jHOxjuXCCOt3dfWouvpxix3KEIyv0HHecvOtZu3UqsabyqyRWmfJnLpnmdniDG6JiynZi+QZ
Ul4jAQVFv5vGxSJpTnlZwvRIyrYXHtXv/mrgP9VQb/0K7URvd2IYIqnoju2dsN1wknG/B9yCsXOI
3yOnsWs7NJyTxGGJa/FpwRSMZHQqFExmkydX8L5VFUEyz6ru7fK9evOwG818XEARcXqHnKXS39+c
JPugPj/sXv6OYRvpPR7x8wDcdxnFT0QsdoxUUVI3OvyMNJNcQaMogUNuUBc04g6Fecm9kjoVCOeN
4YuhyzwLkhD9uw+cIDLV1rMc4oPRlX2V62/FMnqe/iK76TdXh1MTpTL5E7L0/uFz7FYtjkU9ospr
/BfqPL7GWa9lAtOpifu/yRJj0iKAc0sOuILzYG0x7GSatsOXk8a2FIF6GfC2S9UDj64NXiIkIQ6C
NZnSEJLzMVRvYb76dkX8VnFdwuspF50mzg/T20knKoZFc6lrPJ/mUt1L5nGWzJ/fxHEagXPEjflT
1wuIAHKnJn90uliJdhdDT+fSak/sqL3cWfptoJDYl/TDUIGafbjPNDTXga09q0Ebpfes9vJ5zJEc
95qQ8ktul9Q5haXGhK5e8MEpK4lMyaSK0DOE16I+x88HBZuf9GaSy8ZEMeOcjZxekdkqHBqlvn0G
6f3TES3V9WcluaCwBv6F1Bj/Gu5wGBrnHzb52/vfsAml0ovGgaCnKOSa4SkAY8+zf+fkLgT0kx5I
NDpRaHtqk/U7vOejZbYAwJ0RmYQGZ/lJElTUm16uK5SKipHaWCH29Pnhk/Fy0lzyNTLgzfhZRa+X
QJ6/jzigdEoo5v9Gn56vG+N6gopN7KU/fkhRVtG4fv25UyoL000JHPjtUUo3jl9dmD+orkVxS7ib
hJTPxZFLIN2nRJmEk6kTcTV0PK46OqPMUoqIutOf6WxsGY0PYZlmMPp2YdqFnum5agRS/VJvwzAD
7/MiM9trJur6uXZKRs4pIHiyxDIXeS3TKIRbv8iC/UQ48XqIeMKqmjRyUFQgQqDaVZstGm3IQS4C
/HUgTOCnsDE62qO5xUhN2A3d+/u2BszYA1qCyBubv85CKfd5hfdXwPl0u9J+i+jpSfD/GZT3nXbQ
OjgZn7I4othnRnVQk5LdDKlm17EXzol8KT5RqV1IinOAKcufWYE703lgS0UdpbIOCUG7qX0bnZ0u
Qc8amKx6dttFvId+uTeQ5/8z8VWIlEvVnMv/tDMLbyeT8u+NLIWoJneNonwbff+G0ZCVGPefgjpL
K5hgqkkUorTTTTroJXjKC4/dTD6T2jP+gygQpMZPguOoeEu/76zan2oDfV4xqj8J9TRMrQI+L+/g
tG4UPlTgk7ukB2UpJVmSyzeOIlMfQZQpOGopJO4bVEtBkq1+4sArugROuRuDPVv4mc6HE3cfRL3r
CI94QlPP13C+DnifZQtHGgySsE1AgXC0VMTu6z59DXT7UZqrbAvgK1Rb5c7U8w7oUPmzJEQWnLxL
scslb9mi0+NWx66JxmlCZK4zCbR78WSWITukT43ySKEEskP93IeMjW33WqM0lcCK6uOXOXIiCznt
mUPc/YCPbj+mBvt+4IY8khyUCnFNCDN5iE8+lzgzis7QtEO5jAzRRMqPAvaIjt2eBFhI00SJO/pe
fo6Ax5hJjg6v3LI9xO2N0NRZm8IP4JnyoaOvkiuf98n56pP3fWDGyg38UwJ9KO4/F88LJs+zHuVE
cfgHbLkQoiDwSU01Lbuqo4JmpjjW+W1Bncpk7KXmFZmZqVXySrSO4PpigJg7kcAkg5ty012hqhU5
gGyz5DOA7oVtBGEwJJJUXA9alpqtc9kCqvVKGnEsjqw8iiaD4gSdw2Qk+P3J1zbxKnM2kIPY9MZK
QdVRzj/P/+vM2PbL2zVYGD5xVN9scYAR+T3V6nUTvYTZzChQp2zRygBZ/clzc600ftk+SRFv8wxR
UTp2swKMl21vrvvgpi64nf6SSQtpYbmvj/RrOpbQSofrcnaDn9pGzDLsoqLrOit9lsZ6s3BjQMsA
k/JrWZecRFfVBRHboFVuvZCypMmJuvIwL+DBR6C0AlrGAz589t26ZKUQUyGa10vtj2UmTkMjv6x/
eKjklia0UDQJumMS9E7VAZefzoPvX5Of8ADZZ6HP2cTcegWskpTgD70HyxGSuHs8s94xSEC07Cdv
Cy0DplQl5p2aEnM+30g4kDAx0zy09JGzJ86gMmW3eN7xUxAFJErQOhCxVv0AqCve3wPkqFUl/IyZ
1Gag/bARxw+36dEY9VOqcJmRpH+rDiAHD37J6mauEsTnMcOj46csMkSfABMkniNB7gYa85ozCPT7
EJNixA2y0KvdXEe4x4oGpat1prv80kyZaBss+eScy8vz2vuLHeeoQML3k5DnxK/iCPm4DC67i+K7
cnFX3vVLF+sTnHSnmLNYug0U7gSoL5Klqv8bNC7OTaxpaOkg4yXzvduTMI74q8WADSrPFaqpifoE
GKVIsq2qDOokh3ImHnBn7vzOR3zvIJ84KTSc+fWAOHwUGdqQw8ppFO5S1pdyDpXgjh8ApBdtB/9l
qTexc6Ea/qV3KRimgPhkT4A6VK0dILaz7BDziChFzJ7yycReEuhXvdsJfHIWASk8DkMaA08aQI0w
6aU5POoq9KVpdOr4UMVxl4RSZlsNIS7T5eRjb1q3Tp9CPCoVj70KMadxKKZzML3Sn0Ix/XtNqkcX
BTozQpnEa2Q57+Mll3GyfaHumBQVTEN2YGzARk11FN0WllAMS26vYws9jxv+ezGsg00U4WWItAo8
R7k/sVJ4fI/2ilreIDVLvvCJupIXawaWLMAT4xEnmHVJVenqThsz218srhKF867WjiIjcKwgb/KM
XxyYfuIUbSC47Nx10sLbsNuhODb8eh/KlJYkSEJRFJJwLRneqtWZgO1DqUHESF0I69Cv3P/fb/VG
riMrc/Wucd1nrSHQqcEPuHTWkjorOVVsp07nNg4sIA64zpZH2+orJ+YI/884fi7uov11w/2jhYDo
+eGJIIIrr/6DnTrR9wtKlya2wy/vMXD4oXdxHX+V63tkaJk3bKSKQY7oqeqqHeW5hXzGo6qIoZIR
veULnzykcXTRBi3j/CxYPP2hPUo2MLx7bNqPuDB0ei2E7EWe3iPUm35JBgD3ult6f0BGygab14Cu
bfU98NzasoK1igiB+YEmKjAgOh2a0zcbwe4gJDAtFceY9UwdMhiHwazFQz7NeQDxu6QnvtI1WxXp
IBWsxwiZIlYkvxtl8iqgFG4be3LXWFc+/m8zEbFG+k/KtRd/RqbnyVS1ts9cI4ASG7DqdMgV1Gkx
ub9rLuxPSgMWjhUelcDuhFLCctlatCgLghJW/Rf+PCmSjxXtBbat4BS+Up5F6JoexatXJ+rTHg1P
Jx3FG3Z6YsXubPg7VMb+jDlQFMG1MtVS7i7NfZMnokI2JbCRd7SLapfh4n7Fm9VkRl0Zx8n/I6pI
xw7U/ZkLj8RXSYbfqX2xyYiCFwyVf025jo5PZewwN9nJONGWYnAFsiG50ia+8LPZ96r/olzxIT9t
zIhzIxew68wOk9jrg6i3a6l3ppygFabEWsz3SY2SsKfpg874/1ZETrlYyyHkpHGyiTSfjy9gi+AM
WUPy0h1XEXogVNfkxgeYbqt/++aBrFZ2yNuXv/DnVJ1h2g94KEeouF+Jh8gEOmGwt+NB+Ose0Nzw
SvRssJ7ZVZSLLtKcxbJB5Lvmq0BQUNJFkfyJoCQE1FyauHA4pkCCkyw6/UBh5OL5dhwb6WUtZACt
O+NrwQ9utPQpWLIlS+V+r6aWFThepcqsXpmwKyR89GzuRSpL4hgCMUlwVbP61LQIeVWWh4Cn5blF
oqpcCB0QS1nZUqVKOOeVqfUynfnUP2nUfEnnE0zzWdfs9Ewz5MoR9Tc+bs0z7ZfGcTAR7m8i5dnX
EA1UdbadY9TYGvXhBmAFlmTgBcnmjuwfRRCzxaCko2wKlFfEF/hUn742QwokbS037Foi9Wc1tMZi
8stZSO9HFBA3J/+HKkl2cOaSOySfAMU/B3mf/7juukcjLvYVNsb0VBRPvlb1kyZ8i7Yobp+fbthS
O+1TqFjvcYzWLkTKI9siQCofD5z47vLXV/XPhoR10ismT1PcYnljPpZCw1SOjfVleUM6MBz5Tzl7
CYSm3HlIFIRHWCdynVAIMFYPoV0saAHYWiHeDrOXjPXkSgc80Ie2URwFWK9cC5QM/tqfScBbL8L+
qB8IdWVAEzRL/7MoNVBFAt52AT84NQ8Vxch+cxLAwhgOezh0Uc5g8NlIx58fPNDOvwaq6OpkpEgq
xDb1MR/qspYlObd/6b1ra0iPiPqHh4Tj/XVmyB4/NlnXrlSULj7bVOwSK70220TXDMHw+z4YPbgd
SK9sFaE56fOKzfkoeLz+1yOwI26zfhs7ZDyI2CCcIb7Y4xxHOKmI6wOZuP6v83t2cqdE1hJQOQmu
CxkEV5H2yX93bDRfT8IBlNjl5ZgtVRds3js7iDj87UoLamBOtMLpzSvLUMIIQcSf1Pg4T8vfODVp
N+DMhbwL7+J4nNyyMlQpeRD5t+7791HSGSCueotQoTIu6SNI+JPjT0UQFv2L0PB7ePuB0L+B/zfd
7kaC58AyHo3v/ND753m2sv4mnRj5JWjkL2q9g8jdsDBItxATnfQHxPQV4O6l3Pg5WGr/d6u9yHHH
7WMeUjkopAQ8Pto4nDP+gCJ8p5xsE+htzHcUiB8hpNiQ5ve6FWobEWrjbwA/glGuMtXui27U/Czk
d2rmZaBadFw6WPEoZmDAH3HevPUhPiNRr6X+JQ8T5J1wVsCDtJx2wflZiaEzdk9fX8vlq8asDGAR
EVaNYo0BoBXt/pxLi2+ekEEovXAaVLckbS7vpvHoVoWhzfvO2zp+9GY7DqkvR1CRPQfrgLR07W2D
6qumIKtu7qP7R+ZWIIIgrOtrdmdApIGttOCuJcTKqdGFHzjl+uZOaR062XIOGTTc5tyu4WH12vS+
rpNn/ILuKpVqiFUa+PD4dXAYFAGW63BhWoQqihsM4etjZ5cXzC6cHN8p4YEYdmOV6oPnmvRZsghp
vNryXCe87cHUKI9rHLueJlr4PiWn1tN1cw1dvL+LVBJBTuERa1hgIqKq0Cd3m5zeHyV8MWn06S85
BfyAlS62gG1H+q6ei68Rq+0AjxSZlF9CAFMecUQ+l0T6pOV35hX+iqRdqJppi09i3gHlaF6/Wb2T
y74VtStqExeeJEwMYz1r9YRTlac1xlGicdwzLf1ji2xVc4p38glEK03Pwkw1UFXDuMY39O88S5U8
bMpZQv2p9oWMJ1Uypb8pbPA1RpuykO72GTDA+mYg/VeGjlZOTUl2dOCnkUbzJz98nc2zto7metCk
AadlEZmt/kLc6RlmhBXsg1L6BgGfUJyWzOmdfUDQ7PUbs9EhrbatDPJ1Skd0wIrZbb59O1fThwLj
XNhGs+8APJbHcsyF94bSfI5PHIt4X064BDNutplrvCc3FBPl8RTxqGCabpgNe5bjhsf4cKDNRyTm
TILrWdvBtmDOH6d+wWanptrXJpXnmJB0GgX3ni6PC+M7fUr7yaZWPMnAiQ3PCnZUq9wnagx92NNw
9BJgcLP3xn0csX035nXLXtuORXPtw2VmK3h92/OcFAdoo+V8Jcw5KzsWQojnISReci1ljqUf2Qpq
bAM6Kqg0+8XlxNlgH0hCVHTmH+/g9vITXqAHVGbbghoHAxv8RziFVvedQ8QpuCjkiXm8coprJLah
b51Mode3BAgqVUDjFyHAMnnthh1ThTPAOiZ8CDEVsSBs9070/M3Vqu0qF3cRX8BoFpqJoqh1/UwR
TiqkODagz6AV8s7S8oR77sJ1lufo9SzjY8lQUIgVwmR5l2JofwyWyJ+CU0yAOGgdTlE+g6q2loqb
G/OQPkjwobxKSxOfwlam7iVEHV5OsBWOU5Qmvb5dHoTek06W8FvLXEbbpbTkvDpHPjAD1G/vUnTo
GL8v83pn4rWFbb6qbwmAxkLA+2wKXzg6Gc5cpbKzJnV+p0KnKnQ6egkp5VjjsG1BiA+mxyGwwjAC
JRpZbhBGAiNGIHwfa7IXxJn9ZSNBRsf+GQvSEbYDYXUuTVJ7GxUJBwfgBtEkGfnGdH1sFa+Qqjxp
zyDwx2KwMF2mw+lEpN6EEKW9ZFFJhiJEkPor1hhsBJ/Uq37ifQ6QDA+Yx+5DHJUOTE5n7SNkO3Jb
wmVcWZQe9zIXq92/usd7siZ6TB6e9H6xdDIty8jtIc8j5WNaRCFSZcoTY1di4J9wz3dL6uqXZUSn
NThVJG2OSe7VJYRZdkS+AC+7vR9bXjm7GQ3SqZTZRW4EGasI+9ceONyv584akszyTobjPZltH3nj
zfirwOL8jBzfgxMUIBt9dV4g9M0ptc/F3kVsUu3ZHIh36XdOnruozElEbqXbqSL1dfi6S/VxNY1t
jtaE2L/s3v5UKC7xQFI6z5kE6WejzA9Ti19r+1C/gRGSgOz7bmjvdtVsEOLAcXvY9lISluefWNpq
wcp71h5qdnIP5Hp/HRg7aHKL6gvCnWzlA7dw/AIQvn2bKCjZ4mctkia+WnNgyz65a/qw8Lc9iq1L
an+lBQBLqyrDgTesDqYJ3tBy2FNN8vKAjcn6ZMM81CR4AXvXdZiU6HPLvjFWPxXCBdeJduJuqPK0
UQ8qyWbDF36H+8sFh0OB6wy8XQ4P25UnEjdgZrW0JFy8WnWDrwhjZS+sxOekjQLMfAdNm5UEQ3ZU
EVZoqjQxOtf5ipiEgTIB/plDrfaA9ZkAuXqk4S5yz9w3Yn4Aqi2XuncrElv+9XbV4ndZxbdUv1Xf
GqMfOZHhyNupnuXP/1sVpdBGRBoH1U2lujstpbsrPXjfVJwJSZ5Be02S9AWy9kNe2xmEBlS/AkZ3
JFmF3856Fo0TLRC7ys9+VIShOgDzDT7aKOdDaOMyB5iLPT/op/xag+7/1WiN2CH5bS6QBbEatltH
SNIoSnT99XYGEggKSwXSa1+ZXsby422CJb18zm2Px6NFs3Ixz5oV3xmKKqbtuYqJHutNRrV1IL6J
1iXOeXXzexLZQVpiuYlvPc8MNCy0OjHgz+873RspIHG9H3OtUiNGR2c9IwyUqoDZl/h2pqFbbSlj
bf3NC2/EXaNHX0vogZ4GDycOgGWuxANgGIs5fXNGEj1BK58eZ3IdVT8XoS/ic+ChYBa4xBrVU4Ns
TDWO5zd7wrE4H2Xt8i1MzAdv13FVS3BF3yxe/3MFe4EGeLYbb9idyP+MyizlUSfUXGRhWmHRFbry
TyGnTLTCQfVVnB3D4v76yR64rN8ncVfdKrCSz9PhM3g2N9CMy83zZY82Qbkfk878Rq0C/sB8UeAq
f+JUo1iNKz9+z60f+J8qHTGSC8oyyDkU+2Cxwoe7xtZMrNUjOj6oCKL0CO+P0CDk96nOh/sKp07U
J3cFvtNhYCHHJiLzS7fSne7SoY9l2tqllJI4TbREcRvhrvcfeMt7fr9nSops35FsbKaDQkQ2MUZA
YdT3X0RDS+E4YxBKCy3YHsy96EfKwxwdHuMWuj9F4ppkXl+nlk8HpygEfQS2IeQwl1ccCbhaovro
c16Txiw8GqyoJNCVI39mEKDhILSkykbJwwkUewy0PSlx5htmgJ2/HAQ0BP7zRmpeVuYXPRPDrXmt
k2+LjQwX83tBqqDs710s+QkoRg5Pnk3QzPHJ1BAXQmMXy+Tkz074AYzUwmZ4iTQkSrB8TdC1g/dr
bsxrNHfYHb1Hb/hhkjWZw97lsPDeWtRFgoVtcEH/jaEOWgTgtioctvXJjFZdt/QzFSUbmgmbxdgC
2jPcmGgj85GkTjHIl7O62aI2xj0evCpV2uVP6ObJ0KB1fHsH581OntQUaFAOpa3ALD+UNLhbuXp7
bwJ0PT28v2gdf+lHNqordmNBfShPX7NNfCf7IQalmf/MOR7fNItMRlb+UfOAQZJ08h3s8wt/Lx2N
4aKuI5m53n47wQJ7RORbBR0NLIRFg/ButilvlM3f2KotbMvUzT2x+P/g7GQYEMkwv6dPNntoWjCj
1nGYHU4Lf3y1BrMeggYuZ2tizDWOT4DO1lof1IBAM6J6JiqWlbcprNSTsV1sAOLiuIvBtv75arB/
3GH+XKL10KAbudnWA8u1wpbEakTPh6YGUvy0lxHCknzrQacZUF/QC8ZhDyuUoFYVuAhRWqXdvG2z
OjYObknInD2b9uV2rFAJPKxc38+6jIiX4IC9X3ysKvY0n3eHG5hOX0T6moD8JUrMZwR5HCwlf3A0
yVT0U6sPoMYNXOuX4pNleyKpZv86yENcnmrVZkzucTENKpn/abhm0xjwbsP+KIoxBicGQqRPEHOf
rbe/hcMtNTz3nE9ikxn83poX3mpZSwQ+RAfHmbM91z5wkzylSU4L9BjBTpr5Yic0xZFh9TXOQM5q
4RONXFmiYE53BwoPWk1R0xiQ2VpxQOLuugXhQI8oz+dNVH0+W7sUjUREWN0/TqMJZ2DI0fMktwhG
7b/bZlCQY2fpwsXvQAVxZVv7RhWikrBCK/bngl4ZRLMLP9pRow8BKKQbC5Dx8UHdf0aCMBzvSXht
QpgmjxeRTwAI5P5inCV9onMDMDkLOkUEqXJAAywCQ0VurbgbbtNZKWEg+8us0fP1YMeGZXifLXJI
JdRXewRE2zUopUvR4yAIok3x/N0Mb+xCyhtonAlJCbIxz1Rvzgerv9U4l7+0vtinJDugkGjvjgL2
1OEaVcjGzas2FcXfsk/jlpj/Ug1KmFdSTQUp9QLS6Zq94NDN0dMs+zfx9XkN2VTpKtogHyH4haKM
va2cDFnuTRmc313OZ0RA4WIr6JniXdUqaJE0/dYeEh526Sogr5ZMwmvDhZl1YKFEgXwSiswKbIep
IGPfBzfnQEREK7v7wmGvyUNdPADsI1qWEpUKdNGRaUr3fyP0BVDxbi1h5SGkhZQO0TImVvREcU7X
SbWYxwWvN8gNWZH7clYtkNmFCyG7p/4Ugw7gBRWU9FQgJHcAuop56UVjHA6Ofe8ZRuGUJShW2iVl
SWvCLOm2ktaj5CLhdTPNO/znr4KvXhnK+rgtk6uxfScY3tcQIFP0pwaFWixRZ5KO1gHcP4P6DtfI
caubD7w42Fyu22jn1mWraHhj089MtPRhQs/GvPRS0OpIyVmUlFV1P9B1KC6xVBILlmdIPWGB2Bi3
/cH2HFlTq0tTIxDwcTgOt4PjR6P/f9gx2ya+lh7T3EDYfQr672AynudyahPAAwQT+XBFK3slulsM
kwJvamoBH3DJKkAJFY53ChtUBoSGsCy3XK+tJLbF7VpLfGxH3qxrxWSGYJ6JgJ7BRX40jLLzajyA
0+Yyb4vj/swCIVbVzwAe1cdvViuVatgPjtsb4VUXGKna7lntCR0y+3ZJtXtQ2n891wjLBxfwKMqJ
AiH7Zq9fQIODDMGBWaU5+QVuQlBYW1fGWKwjRQXhYkPMjbmu7EaX5yu/kXOt+wmB/bUNluasm/4N
3GA3Y2yTtCu4zu7f6NZFR5fgvyeeoMhIcBtFQcPwVJ/aU+ga333AWmS+WUjuyz/RfifYNcLqGDpk
W0y2QD8honIKoxZJQ0BleF6M3I8sIoA4UBrs3Dt8gwrN61cFOS8dG7mo3nTSbWJbXfV1voVg2EdO
psSG2F3JhCaBpTNdqnnaOXpr5jq1r7kOGfNVil5FPrBumSW5TQnwAyr1BVpdpgK4omIZmu1HV+Jy
XsXovqe95oRR/yz8VnoIE8D+nbnA40ynbxU0hvLBH1OjemZa2wjPBODiQuTGfXigZQ1xMCA/TWgr
iGmfB6sBqjEvRvKAYoGdExoAif8JW1rGMvN1sORY/qjAtnU9AKvSebrgw5EnkkrAes4KnhE8w2Dg
dRrBwSWU0RrtqHo5O/pYLezBtsO1abF6mZzDJNW90seWOGXw1oolZ9BnLiFrhazO00IH7Ayy6flw
UTmB2T90UyfWv2tPCPidpAxod0hgx3LQX6htcSbGo3yRxU7klWlTbd6gQ6Nqsw7Vd4qqsJdscUF+
Zl8/pzgEkbt4sSkbx211XzVbtDPl0KwGPhSILlq+iSdz0Uqj6hJ/DrC4vmSj+W+8a2tLBAN6Wiqh
+wK7kdBVWOukwazMfkgcLrqv+fsZv+Cw0iBRjYY9UUlCStR0xwl+KmhqOuBzgQRELwr6lLV0TaOH
/cWEPgOs3cGlPbjtvZDMwv04tBF0QvrPzuzY1j0ZHHtZ90pPvT07VPGoVjkl2u9u660P1GhgG2sW
TxlgPw7CGydqk1rrC12TD9X+ibcePuCTbwDtFGg14u70/vHdl2h/mqM2djiiloGLwtjr5kbEmSpX
yAnGEiIwI3/xFuIs9I6/ilTR+myK02MRvjhG7X6yWscywLuyXm7+p+3G0HyYFQvSg4XzrOUKry5d
dxq2wVdyXHBTrnVTfjIDgAtZUTs9PPr8+tF6Tt9hOdE9QGEsvtI3SoJPK0Rlf+7Snm4cT4beN9sm
hGoTXDfUpoFIAInxncw2Jgsj5BIGTLNelE9vRpjeV2XBBj3MfW3p3oUPEAjygeh2u1o9ll1W8Wy7
BVKECPtxg8qrCsbqQC9tzBTb8WbNh+BTu8+k2htS5ts1cjp5jejUnRgNkz/ZvunQrHywytmMaoZo
Mqc2PQaDcCKuKoWFz5vVyDkcd/Xickjv5crwpQQuXptuPRkHdusB8mCgYES8VALH62WV+WIjcEdA
c8SkBAP9/s8peID87GYAbdFKOz9E1FR6porw0ULGcJV2UvRpmCN8dlibfB9oZRf4GwxDtz0unzlL
uiBVa4YsVBxgkG+lkV5nm6lW1MtxRa87JJxmrJIPeB9St7YEFfnJ5yn9d64vwrcm3DQWCuEZKFZD
4vE7wXyEbiek2sWy9oIt9kgTpJbdIJdA+UBE+ycx6A3h2HEywQ+B9t2emvaaTHu7R7uM3R8/Pnb0
JBzfyjntQD7Y1xRa2/wV9HpMHoV1/Nwpp4AFCoCqMWCLVckW3W3Fx+x/F9l+b2R1prvDfbI6L3Y0
nCSm1ZRfjEpG8qkFWP6NnbSJSPLniwr2Ps/q+NflVnd4e3N2BrG0eyNpv5FGHjvH4ijI+fIpWsSB
IOJ3qEBNWRh06oAG+wNLb38ND8yVekcpnSvQCpWGlezVJ1lYCEdsfvSEh6d/f9w3s6bGsyBmqD3H
e6ZkPgHRmiLPG7IgXdtJ3xpFRj9Gxgsq7EvDWI5fwn8edB0bHyixWAEJR0xTji6bpa1xNVaNRfQM
/wVKDAB6HCuIz9w4/TiQV/bbopb3cMopIi9E5ZZQBWdo/6MFYUzRKBgRK8B/uGpKKF81vJU9tEqT
HLE/MINhYeVNoaxFnsp0E04mKPiHInQ+9DeUlaFt2FdxpKbQA4ITTvBEMcoS5lVNcxWuISFc+9IJ
LaUUb2qpD8/9IL0HgUwR/ZKIjwevaOePNMG2vuMwiw3iRcUjY7cGVbVqlJ9/3aHLk4wxe2r84axK
mdtBbZVXvqrZ2lV5VCBB/zUNrYR0N9YibEERMaeILiLru2wFLknpAZ1JzV1i/HZitF3QYVmVHNvW
JAt9kE/DdrCFry2D8yfJ87aIvHhjOZw3vCewuS/peya2UX7RXWU2nDgLEb/37x6A1o+hZXU/V40d
7VSjIjvM4sPqfYd3X5TLplF+Qr37Ul7UnBS92es8N9IwfO1JcB1EfGFPJBY/2dVXEGsGsjtViOpo
EdvmqKdCUTyHy8DhGlrQ6Ocd6IzrDs14MJImnv4xPTMnnlFWzGi42lghrmPvApCfbZ2TLzil4GIl
/T8NxAw4wA09kmdzD53bLRGyhYBH+JWiBpC0aD6UeYBTQjI1hn3JgJEAW/Vnlwu9MLbeFtC59t0B
BWVtTzGkJ+F/+7Q7112lowah9u9W6Hg0tfEoFx8xrdPSk67DovKsguv8hQesK6AvMejFz3FmJsaZ
ipQtihcfApaxi3+o3vkJMUy0J9KKHfGYCAWZUFnkZ04+Kk6OyMMv8pLnk0K/9Vyc8f3qNsQ4yOGg
f6Pt0rt+hWwahLVfzvwsxIHeESfHJJN/JvKh5RstGeiS9B1N2nWwSa+aWzC5ZanwEWx3dljMlod9
cNlM4X58idhhqtETTP1xPdS7++AdCw7748peGVmED/qMz3phMhzWCWpq4wiqS9SiqixQHHSuPnV3
vNEhCf7GVYqQ8DmxfCVf05vr21ItpHo2IuaHWFtLc6RrpwFFXGq1AAzOboJ6bQylSP5KCLe0ld8Y
7GGce/L+yDe8xNk2lR6i86iZBjXoJWu2t8Nx57Vrw84HjfEQ2hPlC6JIS81Oe0SuCTa2Yg6oPfCd
ogZ4unbJBVrpfauiUzuTXQTh5GGVnhdxxMBAuUVEp/DCu6e+vb4lKQPHEa8VHOJc/Ijp2RWMHl98
+LQRqlfNERpNwFPr0BTTDYUJVdlx8Z2ESr7yNKnLDio5sEN3igWk/F6Bt0K412AL/obJA5qDpKna
CBBLyp1dr1ViyKfpNqpEJGiGloF4yJw3iyuvqm3kzhAdp+8xylyZNbFrC0h9U6nxxipAwbHbuc/D
6NQz/7QJ3kJd6JdauRIfah4eKLijiQ1TBKvMhHlgU5v71pmX4hheJrKwED08SxVis7c0GCx5vVeo
87/l/kqLwF+poxBS9BXtn+JkaUC1cybEm1mXfJnpNvm6FErgTWXZFw2ELxp4EfeEGoIZmjdW2Oy+
u5s3vEI7Aau6pq3TezoJPtPI1bl3iox1VL17c+Zx2GUkLx3p5FpBGq7lgD/90BYgufSMoj1uwopM
cyTuof+hT/2JfxrHXw7YxlddOFxUcpk6M4MMtdJdWQ8DPWSHuj+/9BlPZqg3j8JFS6ARhGbR9Wol
nRSAvXYPXHR/r4oSslgbIHgiY5X0tnuJIllfrQDFtqD7qG1G1Z1Phj8Mub8JUlEWFbDD2A4QDfUh
fku7t+34bUXj2dt1H/t9sZKi8Z/mipofdJPdH9PGmR5Ax9Ho23iYXzvXOpMqnDMGUfTX8M58ZRNu
vy7DAP8hcpE0/ycxGqxKRejO2pXhjLoSdgGEXU333yoMihvEiCbQGleh2/cQbvJigpL2bmWb/m3s
nK2nP+axEHM3f4GG6G7Gs99U9xHTUDwH9cv+lQoxhPMsj4gr7ZPer8VUXxIyCEXH3IqXzDmPftYb
gX8SOEhTGTO3q2zV5LmVf0l0Z0yqgaKS+w586YQkQoHrpQRcMQCgqVeglH0mwLlSM/v7uxN3Qs1a
unEf7AH/Wiay64xvIybMBeUWoQvVSe8yUmXIl9oTRR5YYiYqKznsykKb3pK6gD7l8I07l2YU3x4W
OBUj9LZOGugd2BBTwEB76x/CN5eoyYS4eauLfVIg1rm5LeBMbQcISxFWtydROoV9yM3o799aMJ7N
0swfzIfYlA1PhOx3+qBIVGZrv0NV8f2/ds8PSozlWv8u18O3Z/Qwg4D1jARCfFRrkn71U2eFMmhg
//nmoMQBICqXEx40xSOU5jEE8T6kfbqkCI1BW4qYqlKTJ0FoFNr/lA7LyB2TG9Nm+zFWa5++weNq
y+kN9B5W4RinDUXtRKVnOsZVwK60CTxGj7L4N/7kiA81zAS+7Jlnj+KL8ubG4B19cxVHI0NJe7DF
lt35rbNLtIdPgBZtQ+bUUGW40WygnaQCiJUbhduujFFIt8EdmqvVilkiQwzh5fQmCpR/ajos8Vd3
z8wC1DkOsnMv/TXKEDkW5YBnFEJAir8LnN7ZTxchKSI0toS8rtgcFlEEF7OwqacB2dg04ZOqcjuD
DzVLbdIppmQfJn1Qrc3ilP9V26/KMal103PFaXHkfhVrD0qwVJO8mKTJbhKBHUKc4q3qHUJtRs01
IWiI65Vaq9VEypnxlnBpXLzjI/8vEQ1GugN6fTqOek4rbiAkfI9dkCVC24l9wIpV2fGDpPzkPAWa
LmMNILPhYr+/DN9AncEko/5pBiZdKkNYqZWnmfcVEm7MIJrL2CoFikslKcX9K2Z7+Wsex5XHa8q9
7B8c7lh2vYd8CqJJd0ayqYVhdEGW4kWnrWW8xKDOE+hf9PfuFTkhGhQFPBr2kqM0EWBHMDI9kFs6
Tqib7jBStB2d8ZqGU98186lj4XkHWW96yaErY4cxO11cgjFGA/bXbD9UZxYPbPn2hqjw52LdDg3J
EgSdsld6ckKDUIAg/QBE4pO5RLr2z4Td3/3v17wXN/47R1rABJTKCbsOQ7uDI6S1hZVNrtcPhGW5
IJKrT25j51n71zUoFkkRCGApZSzErehjnoaXT7F9tdmv/JSrQQjLvtXMUdP/qtQNkPliPxAWBLWx
tJnwC5Qk1pGgHk2SRRet3OFC5dqx/AqjL6W2wxU7Ml5/F4XV8wGRDBLyfJKy4KcpH9pyw4aJ/tgJ
uOzIpK2AlnJyacW1SrjC4j1Hj8uRNQh02LPwWj4n2TdOP4+u9HFrDN9E2X3IR5Nz4KUxPOuDrk7t
GKNmu3HgLe8+isG6EN2YAJHcbIdE69/N0vACQ7/MnZixJ8mrf2hmLY7kp05qcG0vpPd3MDv4josF
nQDm0ndKpaErzzc7fzYy/WmMZfUUVHtdypoiec6FX8KQ7InRL8xL6sSZ0LiEg8aBi1w19E20JVZX
ZNWyjYv+YCX4KXnqEyYLuwReP2D1g+pb6XJj9SmyPoNLnMSzMBkjV10/bZGqFrTKAEOqFJIyPUWZ
uJvy1IPvGb+JF8nsmw4Yv+jt2EaWoFn7IoBsyM2HI3xmkVImoEKkcHeBkHiZd8bz4dlMZkZPsxdP
LQgMgIxzTrgCkMf3CswGi+AkbfN65Gpulq7Ptec02gHTopFVBumi3C0fa9ibvuUZYcVoIs+32lIM
XQUpwV98/T0KN5/iKr+qj1+ivnf94rUk2YfU2UGZPui9cePCWd4+BZ75A8LMqg92mDeBtJZucWP+
dFXTQC9ZU4nITT7WL8xExtlCXaQoWmqRYCYfn9kyd83CB0dij+MrcIduMuvO/fftO8nIJP2sQPMp
jGnuBznvmmxdJ8es1UOYMTjL487k7VIKAaV2kf+zoJ7HItjXrCqyP47OxksjNDFLR1wedpoqyOKy
SQXORlqww4UK3FnItZkkAg3kuELXFWNLjMlMYTk1Zh0UQi1lZ63AL6ZCqBXtbsF0gij3jGCxPwUP
NT+1M0GnCHZX+BM9acuMFM08Dpb+KNFWoen6oO60OzCXB9oIxAo8uf4T6PfkWsi7+B+RTbvt+3TY
ucJJzgI5d93dk+Je2sRdfMBYaeVMMKR8DIfNVPO9Lcj1d1CleDvX61szqiqW29pNsPDpaDRDecct
U+E/xQpvfHYiMWVjTuglvIjgFGMbEXfkzS147i2vn81N87MYh4WD5VtMQ3kFOEuC8K326+W0SjWQ
jS+EnvL5fL5/gvHhLsAJ6hf3LAd95TsvfWowK+xZvLP0uPOmmTnHwojIZIo98N2DP/cqFBgwMHqz
ubvIUUNetWvmRDvl4k40mh2yePwG2BQIZu9Eu1czM/g3GZKTdnP1vzcxW+M3ioN9jddcy/sXAKGL
bsLBM1ZsdjV4GGQA76GFdXUMmgWAOe7vLK8QNYv5k8HB5YOsOF2o13uQlfqqvlNurp94wAmh2lSy
MdDxKXy4VNQqK9Xg7xfctx6U5F/OXneahbX6s+6C28Lewwmw6Ux/BYJYECn4a1eV75mnA8JgzVCh
nMdGyUfCaqV1pZ+T6WyADGMU2/MuF3r+wZ1mEHeQNnAAOVl8G65/nhJxgmHzzBLQlyrQOXSnn1qD
yWtj+aV1sHU4ufLUwkKJabzRX1b2asuGW+stxsfoaXTZva6FY3ugppc8Icc+1hadCUBWq6umeLr+
uk1NuothziEG5eu+IgWfHjrevO7ZmNwlVZMCGVtCmmZDWQqVnTSymXsv6IHG6RYevXqIziXVudEu
4VUCSbKAjzGtoyl/kA3B+Q+4FoxZGZ3wc7o6ObugdjR7mlmMdj1K/cTZ6cAUN/aE7NbMhy6XcG/X
ky1dvYnfkLjguxJ9WNCDGSGgkJlkEx8b5V/V+G2ZVC/cCL88lR5gzPLzLnUTr/RVdno/oZJX5F+s
8ogjgZHmsfVKzSdnLHlLlJA8mvKVCXqe27/mU9JXiZgPHPMo4rkKmvTatyLPouIbPwh4qYFT5D8y
dKIoeEH0BHNuuDYbYJRwCtmFeCKg56bMFc+YnevEl3t8KLuX0HhXJOEvUgCLoIr5cAAlk9CJPLKV
v3YxmbOTjLm1JKHzmEcq+VVaAqmwrzgAL8H8ZjL3vFpgKEdn/j53Aa8dMn8BhnSarL+VKibzAXS3
DtPNyrSE+EvhyigJosx7Jl3UXad5HVstIksqVfpiBRNRAwVexcgL8bOtE5yI3baQNXJlYpcJAbX0
EsBNiUGfhCRrTboDoy1UnETGXDE1SAin4Ot3rVzorviLmnNmWPJANHu+e1zrPGz+Z9kLicsxJzZ0
b4VgLDC+bZTyf1zB2SeYneDOvT1NgXHD4ijeLkHD60hC3dx0JSX79Wl9QXzAx6ghaY8oTp90m8AT
4asVALrGlCx/vr3ndfOuTAcCfTZ/vkBKBV5u16cnIscwQmzXDi3bD2kLBQZapzcDGkW52xc/xNcX
CkqUzeeaQxjalhj0uh1vZW+23P3OwpJDW1QjGoP6jQLoz5LdlU9u4TrCTNgyfz6l4FY0TFpKVYbg
Aic/CW3NspWBDuAnLJFBI/LtPC3LkitsL+IsbI3RnBPq88YFW2wIbJ2mhyyIzzv+d6cI81LlKxE1
XMQRo9ZZ0QlULM/j2hm0bvUsSthhrd4b6Z8pUh+NCzW5Q7pl9z2pNoflhLh9wiu/y74kZgfZ63eO
fiODrCzujI8a3E1OAu02xm+RjbAMbNP/hHsoX5/UQpPVpXWyvOt8HM5PZjeDconel207V20AEVI/
uYq3hduJLT5iG/SKg/qXRPyRgFM1yqk10eupnPw6pLkoIvUIHLVrhXDXcNijxuortE26VZmj88Rb
SJwh6dqO6yCE/lP7td/02pDr2eO7O/GcfDpq5Gs4CHztmhyVt1FTt4u48a5+C0W0xP5D9M39KP5A
Lxj4XBH+8tVVugRcEdyjbaS5pJsozg3kSO1b9phvenIX25uDN6oTZVHiboupjPYoaR8+PJZDr5mr
YL+3RwZDqoxTDBOcx3pxTfEqG4iQlUQeVcwgnUrtHMjEyHhR5rnoUS4AevjzHWljMvFYwUxG7M1D
XdaZwQ139bzybkxkjI72ACdFF0AvJTZ5FnShI6mzDKe84sQUhRKpaxi3sy2UpkAS6SI5FyC4SI3L
Uo/hl4Au+vVuzv4HYR6D2ZeuW7ux7Cj05BOvQVKVOiIMBrZvM5FsYDM/Jo62W2SazSQuLlnuPc/r
2YUl+WUbdYq0MiNSlc3EJkH10fr0sO+bxlQcCM1cBAlUvqSF8s55WUJledx7/wOrce5haPrpVs/i
J2ZfrtuPP9QveIY2qMw2o2TQ+p5T4Pjubvsu7lBlZJiJCZZOxA3/AvpEYxJn6agqE/vQUXVpUe6w
D4oiS9nlBQsE14/3w0X9xHgDMfRVUdsfC0QATbeY5Q/To6l865h3DcoXQIGQcchCLV3THB/Ds4ee
RILq1Jxeadb9e8Z3sbFDDkL4N0+oQPOHKWlyZrLLNhSsA5PBngmyhF2Fs96enDd5cBiPII6us1Zp
2o3JtUKBNICabdGWPUz9zXb5XotApAYWbYFMqpfnENyotntkK9TxxxSoKP70VlxT93dzkp28ll95
np1zpg4g5XU0RmqRbBf7MdJL53uAXYO7Mi58FBw4XBA5p1QkhbzY4Omxga456Vzf4G5ZdJV3wkKs
EbIeM+NSKxajYztvxPi/cNtl0yUFdG0oh7uVUu1kmeLfC1BOa0VY41IaxJ9wk6DLT3u951VOgsQC
Pe8wCfyDZr3iUnFnxgrcb0xw3SK2yLHmLFTWtDdEzPlN6kCAAInfrWURhKNUy2jWqtgELFCP9Uqi
/s8ZyN8/YWv7KW2enK0KR1sQwNCEgBpXzXv79xytCBprssinm8L4gbXUwGictNIzmR4XUrcdPhnG
0gKIn3LjvDIOikmivinCYmGS67JVGtnc8m5hT/4ldrURiP+6xLJWkpEhiSDmnIhZuvsrcKIL9XvF
CITiqEQ18RJ+7XEZwj8aYOR+4uEEI42781oNG8b53UJkiBIVpLGGyCwKdAo0JBdThlW+jkNFuMsM
eE5xz/4xlVcYoQfJWER2K7HjGzlTdx7fybLAVarzSxEULIjFmEC0oxvO4lKaLpjyk63bg5ZJvPI/
tf3z38Ge5+cQKStqv8cGNCa5pV2Z4uPH/z6FmFrgDVwtFP8vddtS+RjHYEkpJC7h6QAgh28u7JpA
FQP7RJaLOfbq1RZ1K+u1jKZsML00/EFb8HouO6ji7dR3gKYD37MSrYeqw7+EWKPLvt5mkKU23YJU
I50dAb79E04PuL9j2Vg5Bwb06/PwaTnI+EU+xpXuqaBX49XOjF4NaY4RRA/cLgOIOiZGkHpW9F/Z
61JqAM5dNxgfqqiGFSSNKI0gTxa2spGp+l2++KavVIotN5CyYzTVFV6nGZ5tOKA0ADHFP0JJBU1e
WwztWO3hNbnK1on4qGSNCwcgPu43QM/+EjnHtg4s5lZz8wQv/pbNPss7pfCulY1rGWeyrerH8t9r
BJNaxTL7lEc0Pi6UlUfrrJ5LdNY/SwOv5c9E7l/knqF2NsjaSBIoL4cAbiWL8DsgDmxtJQ0oInhr
hwVGkUf5i+yd2/cRRu2+sUHetIUNafNE+dB7teACYeMe2pZSwIqzK51illiCQTSNKfeWwmOsa+NY
GMi1A6Ia8UFI01oZaFnnLZuG3vvlxKo36C9Xbm+xTgQtLvdtv70bZMhpZBJkGu63jeBpIHrEdyed
lSB2k0QS8CWjRH5jCHb9+XnjFCgTMCXcQxXTUffSP/EgNpvP+fTrdSIMj8Q+YtAp/UU2OMZTft3z
s8NOigyIVYIfKfN7VDDBAsw2NmJHYO+3t8yxJB+RhXdqoXViJ4XkGesqFzjWIv8x9j+cteotJjEd
1ihmZzQ7df5AE+b/Ys8rsIBBN851yZDW3kiVCw/RE+PUcrrXrnJ+Gq+BVmgH12qeTReWZX51GAmO
cGnQYGpSKfkzIewoY36VELpveZyIpBG9b6URUXwKjeMqulgOp3TmSc+8YC+2sAVcR6pSDNGyorFu
RCwC+Bf7d9JXSa++McBp1GWWwvzUWXTqAgStXj8rKwDrGadqGOLDrTHA1h031Ta2NjtwxEtMnw9j
3zUgFO0JpZN18Rl54ZKC3BEj4LBJDOrrrDSQoN7I2GKP+7OBoiN4IOczUVArI82p0/J9CryBxftJ
uMaTK6Ivss/otxcaFUlpk2ZmwigD+JOduRZbqaRIPk39Wdp3vv3gqSNNF8tcsGsUwQHhPpSicU+3
zAicoArzCfxYvpZ+BxRsiDDJS/eQCAnvr8vPAz26ofdT1M70t9aLgwG87eUGy/S6V8T2h60ypoIT
vDi5psi7z2sgEHdMeel4Dmep2y1qYo1lsQv3aNOyuP/8v1r939Ka2/L1uz/BvSUIgs+DLUgNgIJg
GF7EXRGogFvEBQkQNoHYMLHqQhgCj6sLn+qo9j9UKZwO6UQ1WE9Chl8wR2m7UlQGxg7XITuh127i
VHsrnzBSXqT+kgP/gVT/cpkGVQZx5fezcGTjpiTCYvmAfA63iNS+SMon2/iolup1yn5vcC+HzumQ
T763LRGKrSNbWBn2e2rLHzLJnJmNke5NTjQe7i2orh0lNn92oGPYpna/gziTtpa0YmHYp6n8JKoB
9f2AMrsiAI7smSMXmp2CSCUaK0fzPmhrsdO8YLmG+srEjdm4KQ7eZhYiEIkT18uu1wSpCQRM3hnD
8YwnxMatXAog5zOtaGwzs5DCCcqjVE0NV4/E4Mrd/zvRk51JS5UEZsWd+isf99SfoxUcCldmcQuW
4Pc2kdLOgV0GjIGyS5PaA4TeETA4bi3lkDDmCHYLoxtmE/+m+lFL/rKsPQjuVtRlNp+Y5IdTDA0d
zhq2/kZBmQzMhFix92m83WXVQ/kw+ebsuMM7bqY5CaBuK9d2l0U52dluz9WS37vSx9MV40Bz4tHx
+mt5sNvzDVYBnBkl9eCzCrxudkxjtrmQtJMxsiYUT3LpXaC3V0daAwsk969AvzbnoY2LfqFGrkrJ
OTjkP6gScq21tWu73vv3OI1aTXNaus8QYR7cRJnKvK8RRNYMU/cGLjI7lj3/NaV35iW4IDaZ4nLa
/cP0l2SkS5m/UNtaEaSMtxCkO4fdYqNub4BUgpNQ7AyGVpKccLh2lR6oUbDXSCnTgcMIbjJED1oq
AUlsqZfqK36qLDvEHPsj6WxRUYBudg6xY98WgvtOib0sUiUCC/MgJDjC8EFfCod/Nh2v1QahuNkn
hANkDVdPC4l0y1D+0EM7snmCDMGHm1JDL9N5IntIjFF9xZRk7Jocd+hRxOLa2vVmYOEa/ACEHIo9
XF1ESh9WQdwpTJ4UNP0Q3EJR8C6Cq2lA+BYQbNEp14cMXSWwDxGCDiFBdGxKKSdqkMrSDvMHamkV
hyRaBFri0jGVhaXot+QIhtMfqI9YzoXTlh2jJ1hslZDMIGUpP9KTnIBE0be3sMHRdpxsNrFh4Y5i
ydcTn0J+GkzPuR+2YR4QinsUSM8/FZIEd4HMkhYi4m/MZfOQ3CSO663aOPTMotD/BsOS9yarZwFJ
Keuy/6saq8kxZPkIYCBEMrQBPUSBNuS0HN6Hr4jfwcklsshpA93f6huzIA3SpZRg0fufWuE6dK6a
uvAcmTIqVzeJPx4QkNkehOQND1RAg7iP7KYM5ZSNmj3fU0XoIu7q6b8hf/XV/dpEJ2NbwxWG8D7j
cNB8FIj5Vu8xKXv2mvfXoiI3H9RbzY5qaK1AJAb9/UdMiqXMMQmw6u4zepYch4Cu+eU/7Ksy+SbH
q20ePhX22w1xGsxcCV19Pl1iJKFlEJ0PC48YN0BTb+xnEKznWzXQZTsD8mHO6ndxckkyUi4Xj/kt
lQC4grgz2cMUChouSzYX/HfK9j3BiH375A4PX/e2bpJU8ACSBClgsYeaf2pCCTY6Om2dCJQTtvy2
EXNErAXrYuBZkZsQXNA+9G5ZwjwwiDVgNGXoHEal44LFUFzYxJ6tnqnT5IjFqq/GV0iHHyeXfCTm
5q3/1eWE5soYiUmzOhV35coCmWLzjSCLO6NQq+q0BzcVKgcFX3DgXsL/7YBjiSL2UfVqvmlTG3XA
K4jll9YSOz5ZtJYLdUtxOqDzo/h/5N7cFIIKOApKGpg5ZCrdP6ep+Zkpo5CEZCV8EM0NGi5S7xjZ
Y8S/3qWsMwYS+QpviXjoczgotOHi/LB37Gxl+pGllbuX5bU+81B2x0b0CTTIYXa/srkaGARAjdhr
uZPS9Zh8/4JmdS60JgflzGaZSA315VyaxNBE+r2qYcWcLxYR7RIV1U4yydwJd8N7qJGpgly1R8Gw
T9VWOm93P5/SvvvwW0xBJHSMXGPE6An9RsuGk3G0iwCMqiSXVxgcT1GthheL9rUJUrdilWW4j1WX
oU9ZWh0H2FrbipXI9IdOMGI3D4zlT7sKbat9VVVYkj6R+8WvdGpPcgKrkESi0GMfWfYi7lrGI6Cu
USWR9RrTlBZv9NNkNqnu0g8bL3ngSRMNmWLToFcMKfuDCQiQHGdw7SZfAbxFZHS+NXGb5nkO2zIP
ApkFJe+9YzhHeVcyr/2E+p+l9/UMuqCko9kI1gGzsjxkjrd9GF+iY+/p/eQL4GXoy9oxwDDOtUCy
Q6SS/FnlwShTp9env+UiwuYA61g/7xFF81NBcN8/h54kZ++eYUEzxi2RqDqdV7tqR5O9innAq+Zy
zskBS14oL8I923yuvPwX2cGhHZTdtBdF33lvuhHEY16dlY1akw8MzVFTzjsxl3y2KQnbs3knXM+x
L2e6pqpAVvzjsnbgzhvV5F7+SxBvdtUq0U8S5u9ZNaHgpg3p+CSbMe7+//UUm1Mln4DlXZ6AAjPC
ntTTbC1amSjN/H/FQhx6Bg8o6eanD11dtZ/WFVBXY7DfELCTiR7p8CNVXgdzwpgorO3RiyP9Wm2r
S3hFVJ6rbht4cmV8lWU4oHJ2nV4ahlK940WPdDHP3J+3Kg+yozfrLGLkWNqA+CKtpMXH1znrcJvp
zpVbAc3C3A1CJHX7Ou+qtSbBSMI8N3kUDOPc95mb8R8j8q4jeeP1SesfuYha5gCrR+8TKfXZBinq
tmHULjkDL3/UtfAiVfzdeIjetpgMzh5MmMxwwfL/UY8vP2h7ry58n0EeryDT1YUGgQn6lUTKuUvv
vq9lOSOGclvpiAdEUtfkErir/TPOTBbnmNg/7h0NTX6WIRLa2fmVimJOgThxxIERCDgaQGiUhwjZ
zYnSjRMZoK13wW3jjINDV+XCLXaJOzpnA+2ttdsgyRZ1fP+8YFQv8XlMCvhQbzF9lfY9dNmhzBSw
DMUT3k+Pu5+8yoX07+yHXVryamoy0wI3N56/N0L7zKtygz/E+gKy2SMZVIZGZpqJr6LifDDx1tvy
ll5tm+Bp3axCjz4WcfSAJiMsyMLwH+ac2irDmXrxxqvrbw68RVdjjhfu0k1YV4opNIRHWQ/rf1po
JCyH0XGNcNcEGSrVXpE4OO/gyHRD3UsLt8TNp27luVISxucUdyVQ2Q6MJfYNGYN/7V7wfFaTpsQ/
xfREDNWHgLxteAnqd/h3HVn5YG6V1jgZ8d9fLmsTV6sYRpBQVIw5EFSEVYN75a1v4AXopyA9tCzD
J5pzHyW0/koPhwy8qKo+Ld0JMFE6HVkUz9WcQAOjcfoMECCCRpvERC1HAMyM6k00k+u1QxMo0J7g
/RtUosy7L535y2SKzHXHbsFhMUBpqoWCLiR2sSSHf9mhCOsKlf4iNtfWfZAejwbq46dgIwezhJd7
pqzRPyrbABuOYvHcdoJim7NLgpq3qfnSKVwqQ/KVHxOVdyCtUMaxEj/atgNXulkstVKzoKbvPIeF
z/7Cv7sL90d4TMTDh9A8QnwS3ttrWYuGV3W+gMKoDTTDcLMxWIBp23LDl148OFyp/ZeSeyVTskW4
xaWviejr5Al3F2huxTdoNGL30u3IHRwlqGq5VJA4j6bJmWLdHenlOKggaTLHiul4C6RgtNxVjBW1
foaAJtoSIGJ2s1Q+XSBOTw8MgJTzBPP1evWn0L8zBPotJz3mkclmD4ffg3KymIxunl+XY1DsijrO
kHpjn3ZF9e6+vnBiaCCHJUzSu9ksD8yi/DF6/qXE6OfRYmSKnKCbWiJ4fgBJtDTxkakBD34rn8O4
X5Q5jw7PA9xso5xA4mgLdCKFYt4z0o0lyTfHKe6MpsMuuwGbyzvIGaxyRI9du/Sivtkc3O2nnnOd
f0FxKb4DM3GiDvQhxPGtwLCZQOdyZ1sLK5wwn62jiQWcynqVS3O49fYspWtkBBAZwAPmg7/yMO6Q
5X21aLq3YYgvpSwgB9hvkCHVgRvnJ/GE51hGCdTpe2X9rA5NhQyx5R/P/hfeQDrDvn2G+Qjl4JRq
P1RM76qDTwWRCTX+di1UfqoJ6B/APILEgwDPVCmb11FxR8HeVlJYe6RlSe/3O3bRB0Tjca6/6CdV
ya5U2UGFtGw1VYhx9N5L41TeAuhx+lMo5+KAsUnDGZLkQAuY1ScxPHw+MO5//4LL5/7YORnP1QTx
KTUp2qy/4knz1CE3MnozXFeqq7QOr+wSisKg1cZp4U62cmsL2UaSL+swQhc/+xZxhzxLdr0eCrXW
aXVLEDU0pD45FwvyWM6OpjcaWr66+ulEJkp6hOpelhKQ+gL8jjh/b9PvFq0PjEFa5Gu2EPLxs5+r
T+HNLYO0T4xXaSf5pBE7N3LCmKUtRfY8P795FjY4LFx18YICHbypF1QVAa0PuN3Lg78TWvCzD6gs
FEyn5zVEctWuhPyj4cVT4hZEC7z3bl0GT0Qa9LPDz1WjdVmDVgFTEu+vO1Rqbn2JsSbA+E09anJ4
as1y+AWIdPIPGxiooacKL/5tzWYYFagfWtiOlgHeIERGLMBv5t0NIwYK6FEC2G1wIvYWphP0iTT/
3WmyWyWSQSvaWwajgqaVhQM9uAcLntDprMqJppLYeQjhLKi4VQJ01fpye3v4N/WiCYgmVKk5AG/x
Q0EjHT+3+F2yYh5tIXIYcFo+xYp/oz86X8Ea8qww3c5ZY0kdCMNXuQkh8XYK7+iUOQVmMbRQ31Bt
Gh0g09zG21YUeqhgj9jyv1hbUfj8ddEC4LxGLjsG4H6OfGB3IMlcDygBEgelP1YBOJdbD1jx2Smh
TFjYEYvwFx+ZRv+Av/nSH1eG9SiwMShbUvTfA2uZBheJ+lM0AfwUL2zMrpwaUAGGAwvmXCGr3LSf
PnJO0uv2uq3nLRKDgaeMgfNHb1H563HgVyp3RGNE60wQYS+u2vyQLOekSkEU8CyvSUltbpv1R/nj
RN/9yxIvI1Kf1JGGQvfnSvL8RVdD+oNFcRmgBNrrctSymACdfffYsLb3DufdYQn0pnMfe5juoBLa
jE+OxRlohwguTQ2JklaGXcGRPwV+3/9L0ljVZT3g/ijnPNk6Ua0LqQI3+UUGlDBaqTjDjjN4nTXi
I2y1GSv/1YfjrReyoyqsmwNSBJGDVu27koV3nfBlVJ2gXLqcqzgk2hfuhu0XBqtF4i4t+XLNiAZZ
166EAQrT8jNAIYCqYTqKOIw5JY+WbXoMYHenUDs6y+cKGOEu0lNiSmkHgYgDd3rNC4ge2N0ysX/Y
hm2+TCjeBJMCgDj6Fx7X1dFgqnR54Y+Z7bopZvcxoQUiaVQwDRssw6ZHLF807eNaaCG4lVFx+tTt
B+tF1ojgeA0kO81QyP34ey6Cd+fzJlmBJu3zbzAlNdZM5FODXUVpYyM3VTLkY/+Iyt7UWJWBgRmW
plQujpir8jQ911Sj0IEb9nhCD3NFosH/vurgV8GKmAvLrwm0mgX2F+baeYh9PzyhqKyC+wxY/j7D
McaYLK9QKU3PGPCZaeUT7qmHS0fwB36PsengrzbiS2l0Zi1jqgpCY3EkfemGPvHc2bMQZ2zw9Gip
Od9Pk3mTVz3paKUMJj2NjU4deve6r/Wnk8jpJ9niMoV6cy3bhtk6WZHOyE9naJ6GzM7dUkhkKRCI
DtxTpTAbZntv3ygNZ6wbpJzrUaBCj+kNDRbvKoxkNseJ3htli5fwLlKqzVK59eY1WOKBf70I9w6+
3i58gwEzHYL9mablIvg3WUqL5HYcOKnAQPr0IB1V8+NX/CE5qnDEmou5q43IWG2RuUbcucUwrwuL
oKTN7GSTakb3A0jIuGjN0uDiFynYCyxUDIcPPI0+yZWwWH337VI9rSo7GfLeJ8AWriuewZjT2pCC
Hre+ZdhHiDdS5n8ZBQqeQv6eRS2bIRyjbqFJIzlW5g/b8Zrvf44Za/EZTyrUnUrSwcrWMhrYpC+U
RkQKj1bXpXwh6PkFxHXiHxCNSH2T56zlQkFtznml5nZng4Z8t/IeIyqjtMyhM8Sf8i8RLVQ/F4nh
Q9xKjfEYApCXgqZAlL/+66xCJLWKTp6nyIxdDV+u3o2Hb/Xe4fvrwD3dkwHhEBUwXgNIKl7VG+4J
Mu9hNEUx/ohg2OnPLINL6H7BPIrQIXqBZt9BEBWJhC0epdqJYak90PHGjgZmxBkQD2Ha+qDGkuAM
jD1XwpVfbu/q3KJNDe7yN/X6UfxtkQ+sgVtB9xcTtee7PiGhBEBQkkbSYkxzWimXCKRhXPvCAr+0
gvRlv0ooCQbMD/bCFdawBG9cTUxpFC4jcPVBxF+DKBOZZgWuDg2uMjEEP6UzHlICZ97okzmUDfmh
fzby7ZG+/s99yP1a7IRLNr5qevpO2u7sBm1LHiF8BpL5hIzCXvb7/zdpVt2/oZPhysUEIAyMWNbG
NF3t8N0TsFBvYlBkkabQ7u04CVgDpnApXZaJLKlbHPv+qS7TwYw1hjvsYmlpIA7QesIH6ITWCzgL
KQ3oAmWTakTMbky3Spgy0deWAtfuWAELD6DJ6yBIQHRa8nqPdpq82CUX9gLMhGv0KSlvXfd79595
jiAKXCH8sozkxlWZdmXllfLdnMZHr3C4zpeOMtdgjz5q0Vb0py9NPQjTZfnQ3k3Kbp4wJaCO8yvc
Ppo31Pgw1/xk4ENih9hN+qtapOgnsbZW+i/Ik/M4VKbCeP6xf34ex2ZsSKtfxO/6rgShs1ZUnyWF
boNM/xhms2DoOJnt5YxWi05pHsF520qW4Pl8aaVhOeG7YR+M8tDjwUhJ8VQBBq62Feyn3GYCEgD8
C2uLkiOKRlOk2GIs/aiVEZuWXgfQBTGsMusgc1MvUu9bu4uBNAvcPM07OUjSDJA4KIhITlzA+thu
RpYRgnStspD7FJh6mNElJnLkXK5i60OmcloVDyJvAfu41NDtrdPqyXZSZC/MHj+tv8bAXJvMPnNa
9BgpH8wP4BqXmN2sbqRpo7xnvtVcbrxBpzuw3+56OVt8pYbS4BEiIsrugORnnu3Sl85Wx6OxpWwR
cvvJD8uMZ9FsSn9I2l5i0J3IahwDA+dtVBUxV4WNkVw11QCZcbWw4mPfKOQBcW4uLYrRzaMPDQ9r
SLNu9h3bQ1sVGgCB8/jTACrwNc4EMgkIa0sLjg/lwGMKwuNPbMijYj6gbquj+Yn47K3/EVMYBpae
2fKDxVEx6RPAhEKlzCkNblpJOkuNctV35uROI4YnoEWuidnyuTluncc9wdxMXhEBH0P5mnk/+QJm
BsdIQtl2q3YJd5C8wIOrMeMu0byOtFSntDGv3Wadg441v2uKm624iRuAyCBp3VrtzvY/YnAPcfXX
6RUB+jMhu1pbILM8q0asFrHnodfstekr5OhuW0Evx5KF9VGhnBtdIZyNWe9uhw+KTZmH86g4KyPj
il59XlzjZwDTEq/KEua1q6XVUhfypiydnqXb1XDMrl6zRT0P/g4DPzTM17fkK89RVL9CFriOwmOK
6pH2MYxvjkWnEfp8Mx+JWb/YspguZ6PAuQ5vKMeLkwl/jQOFGVT3PnNZVTb7g5baU2vNYFsZAqtI
Mbpy/fm8ZUoGsnLVP/6kiOw0LSoz52XXw1WFyLu8h+LJm1GK7B0ghJ4KGLamYxOVYDEjw5TeEqhC
qEzs4j94Zf1cvgzrxEOjgLN2v5YvnWpaZW580ytMxTRaRW0hms92Xoki/9hs3r8fNEHOJ1JcKxT9
USVEzmX3oQbUbCsLNiJQOuQKmU3pbi/P8DprUAEPyOLxtJMQH59D/cAlYwTs8jexGtcPeF42hUCV
fODSBCwTss+yQ2gATTXuCybtPRiEP5cB6TXvjbE4ZUOYfBFMF3Oq74uVhnCi0ZT3zeFZX+j2SfJJ
2ZwJFuRB/4jZ4gf+GcGG/MrfOeFxHHqQ9XjF2OQ66wq2tLm+ctV1gt7xjic1N6YAhNlM3xy7c5sT
FYl3GXy+EBPvWqZ9Kxu9zfR7mWbPTIgU+veYc+JUk27Uo9MXioEf65cWy8HxnRNaaAW6/WuHdJa1
Ikag8xeFKFx6FZeEYpn0cNSSchQEMmGm2IxpvDRlV76jKIf3OsTBBBvTQhW1CSAvFN4BCBndsgyS
L0+cdYSP0qisXUY4yg9OniRuv4dE7v1dOaD8tbXwMNJxDnJ+KUl/HLHqCT2p7Cgy40Y6jJaT+dby
02WNlqmVlqsy/crb0kwPS/Wk88tiZzcY2bYHDD80NhtWJy6hcDkQk/E9j76MPfN9e5w9Qer/SuLt
t6R4hzFc4QzMObgAFv0IXuXeintHwnHnT9Je7ixnGV8T2MoRpDOo3Qxu2Y7m2s3lnExjAD7nVLHN
8uoZQacVV/qNsk5qCAL5Dnqv2dTc0T3ATlsSpKSMTpaHOEQJxd7mhllATAyidPfu97jJRKxRgR9o
o3VgEx1PNrzkPuPi5MYA13hPwMeWrc+MvHfbAhdWPjUOBC7UFu0XGSzbZYY8ndWH3OJumcgoIlpY
OxWJatIzMLxBIzNtFUCx0PG3eKkJX9q1Y97HUOuFeWoveLnmmwLwA/ci1JDLLKWSM33eJwz7tzua
H20fBTh7KSEqoCdiCcTUxmUOOvL8MrrPpON02bOzLv/hzTQyTpI/HoVUbJhEz1X8SEIoCvXfcYWs
LVBz5JIwT7MmYbMvcHze2W4yVnK/VIYIUNs5HLbPO7qJcKevX4LcoGdBOBibUnhim7ka+Pm8/xAM
4f7USXhMawESf7R99W40enOwauQjptKb5dax7cvmhN06DaJ3ttvpOCt8O+Uw7ffJV2lB34YJFd4k
dY1tupOk16TH58UPIoR0iU1I79vpDDa7A4wGxgnKQAly6ZmxVjKnIwEzHCNIkMgvuxYpAcM73DMM
EPAuXaKOfApIEUpp2VR+eiemmqBqOftrAvo0StoytXRpLu55YKj6wfKmPjTGuHBk64CPzvVX48/k
uWXkR8CM6oDzGCYtqMaxUPkYY5AR519jFWlD6iMHZXB+8ZvlblxDALoSKMLgmebidMDFFUmTbwx2
8BhLYC5pJnQAYGoRWFc6dA+3TQN+JZj3Pv/nMC8bBe+4So+vFEuKtnwtp1j//BrqtdzU6xCFk8TB
YaWz7q24sEaUj2euAmKY9wM5fW5ug2tTBocWvJkwV3+PWm5R5B2wDpKfsMMhHbW10CSGOIJSUhXn
WduFJBRV5uDtHzxq5z+aSagfr5ZgE9xL3PuTSsVbFQ19x7PpU1hVLDwObOZnKwY/DpWA0WYiIWuw
Ywnxde/4pQOknI/Ctx1DYmf2T3C3AjOGl4pfB0FSrQu58Hvxolc5YJvbg1CLkpCkBcf2pXa2Bk8o
QRHzpgbhZPTIeFZQt3ORdst0Xnlp7N/WNBlQnBQwPRxs59y3mY0YnJlj0Wx5dIfORgGB95JXAvvH
BHQR0EUJ3+Ix/5IHUwkGvvRIBckGMTdF76cigW8hp2me1hlPQyDgytXGac5pJMCkVuAmQCE5W5gd
92zwanih1RUnpY9kaIRnC+mB5XRTAVQzZBY7OS9Hp5SYnPCyrlM27SZ5h/4MopsOmhSpReLuuLYx
A+hohJmJvgQouUc6cqZmuenY1B7JW6v8yhsuMWFrejNg6QRoMs4RnvO3lh4s1d2V9axdFRk4BdB+
Mf24VfyXdJAAshahlvyxYcVDozQ4NxwYvylY4PN+enVijw3DJGnL/qF/MuLKTN2q9c3xGXHDaQ+H
8AUZAKVUmPk9WeZB4UJ6p477eWN8aZyytuGy1BMs4pOXKdS7e00H7w/vAm9BjYV3KEk1HiFFwhDK
MUCYXKB0D9x7/ZwVTZIykIlOEs1tEBM2jTX2bsZ7N/X8fKLE+ZZDaV/nmmwMuGpB1R7+FgzpTz6l
vUWDNCR9ph1/6dX8xUG87hvo63S4wxPFebvf12NsCbkppyI5hVDT5VDxR+d5t1PoO5IZojkWnHLH
+2e4MR3/Cp/E+vEpwf4JdSEU7f33EKdvE5g7nV1wUwXO71Ms6oiglwxw617SoGBSPEFR8UCN5siG
I1IoxAViti6eoxYYkJUMijxvKNP8myB9wk50NPhJuEomHRBWS8bTUwqX+T0ZwpGKc8jnftm/vPxS
8bsVdOhyFwhVnyFHIr/WnyhhIlOw0rHi4v49y27A+RxP1V8igf1Rx4WXh3i2o+vKPQsjbaJBk2Yx
ZGoJhKTypNMBEjKhJyhknHDv1Gtkz80gjK/ZKcDh5Cg0ItWCewI8bTZb5ADxjrTAfkq4L9Rq6lfD
xian1R1MFo8dliKacr4GLbb49+opY0MEAsZUrDCKPEVkDJsHx75vjq4BaJt+FjblDCgbhYdD9Pfd
ctsa4MPpnfboJTwU3Qx+P6C+nZ5PBdvJ2AtxZ38+aO5Ax6s+476RcRfahRlZJSGbX9onFVLnY1vg
RD9gGTa/o37byzcCyCcIzgYp1CMp4a+HdwtoA3o0q1IL6Kf41g4BTjQbjW9LiMXwkmuEwh5yb9XT
F/KeSiJUbUWdNQSGg3XCQiyTzHKuUIBuevCuC1tBDRXgJIB1XgdOxh+KbOBzZyVg4fi6S0y5Rz6r
nAkJQRH76DOpRYSsk78V8l3m/h9r0aEGOvpDP5MK5H87fZRQ0We1gb6af4KR35b4owv2MjCRKbn8
UEx76/OOxt19uhaIguTmf7Mn5lTzkx/TuIIEQOLbTRQ9KWIx757SuRCdVakMzWY9nqNIvahX/ZZm
M5QMJRYATBf8y9YEIrTlB+exNkddaP9wvFL7tS/ijOJXzJp7oUKTqK4T9OaOTosy7/yqFIA0g5mk
MKpQr8vi6z2HOD3lcEr9RrsMLrpGcXgW0Eqng3oaDzAxskBXHr5GauWdjI1BPxZ0Vj7VGW3YTAms
PzfNhDm8VbDcTfg1+fMbYV7c78XOlFJGB77O/IOKy2IM5mMWZ1D6shU1dMhHXlwRK2oolmR4o8Rp
whrxSMbqt5vWl6zyCiKGTwLh+QcGfOpJVDRmP2anV6Y5bO8r/sT16ARsNt4F7UBezFsGiiAiN0J+
aUZmXxqyM++FRclxcuopFgAS0tzWQeC4+/Jb9q7/TKYUNeVYvUSMvV8mCo4H+QwMuxWN33+ntyzp
A6AilL+KEfyV8UYDYaxMTiu7OsJ00xKgFn+VozAzpc2fHYtaFI4FZFeDo9nyo+2XbswbA4Tz3z8y
tF2Jpqawtrq7UEMK6rs0FALPc4AifA0MIHk+XMA7My31v6HbyuUS6+6BLnf/scrgUkIk8ED+XGzK
o5dNjm5D6dK1v8wsRabtg83xvZNUEzw9V4fB4rkjuXghBqgv0MqHJgLDqhI08tMK+/L8sozwcw8O
9qdl4f7o5A/1xWZbfabBIGSOGrBElbQshNNK0/0u3pdx6CAEfylI3RCKw10ju7JLqhyrxYdGfumw
ugBjAo4ro0O7t5r47oQvZ7ra44Q+s5z2lSdYAHprbhoyf4LCTFE5oc2IbirYNnsIUGQcnVgS2ILF
niZJYSqOcSjO4i1Gj+9JPb9p9QmlnTvaOmu4hMhYnLUNf2WgVUWB90sMcgjaPAlW/0RO60aA2//Y
g/qOlk8fQmBkW1MX9cs1Wt1jt/M5uLBLmKo80AnIDuWkOmoC/UDUDJmMjgAUakPOBW6RiX5Khdni
PAM48+bPXikOIKwWK+zqzrvrS8sfMfmRZtKIfxmlvV4j7i2SWbxbcZErT+PlGKijoZ8OCtjCnMpj
DL2uqRq0r7QEt8H6Or03UNh2fXAs8vAicjnrf3ra8YBAxiK9236Oe9FbKZNBIGAiSUfwrKQiLv2T
rxi2Z/YD/RPSqijproZas4ehQ2D3JuvtQyYCDnYl0BL08sngYmSvYsEB6rMSkJmd14J+jdooVnaX
4hX4EX8UXTY7yid2FNWcOcEz6HUM49zNIMLFShcKBZ0+D7MLx+cqYoHGTZgfUjxXoARSWfGjRHCL
2RqN3OG0LKSHrOnTWWir78tnYux6xm5Hap4S71LSzCWE5KyzW6q+RvbPa2CksmBrHjcysdGUPR/Y
EghFSDQXwu4UEI26bZWTEeDVnGmRcVvXhgZJfpK1EQ4kBsUTxS27uwce5wUZLo8BKwgGLm9KvKuz
U/vJqF8roFR913gxLIU1oRbNlX0cNolkLLDWEN8qYyFL73r3G005p11nQYSpxY/kAiYTEoSqNKjX
CjKLksNkbqG91pUOgDXYDCWc2EnO0bS2lpd+Rtj4ns/Mp1UDrvsYZu5Gj6lfDPVlLrNsf81zHJGJ
c5Jv9r90ASqDv3NTjWhx6h0DyMg0jQsTLs2AfIgjDV/Q0bb1ArSzUplhI+zAQWqKJz9am4/gbssi
WddupuGhcLo+lu3M2uU7cMTkYSGtg98bb47lzsGauxn7KKQ/L6YsSkpkQSMghmonCR53whye96IM
AMR0HfKmNmeBH0VjhQf+HSiLj9zQe23OACyRsMKhhI6w/G5uR14SBNlhRe3wUaGGCzNe5xOK423j
uZ4INqd+H5enZkPPt/IwDkGhenm/HEvx9lS7K/OA83pTPM8KavqprG7rxBj58F2qKZ4UA1cgUjiv
hC4+SsIhYglxb7WYosyqaLrQb/CYzpIgGTLHjL2iGDI9g+eG8MWEz/r2ufTsAVAx7wezD2HlUGh5
1cZNlACKKLGTHVjrnDQCyjtPPRzlJ6Awczkwv+jzxlDzpvInRvJWlbqAE48QRXRYORANNgOm40CE
GSXW1b3JDLKfXewDDNEEzG4OTHU4wYGCB+2i1Ny71LeB2efbJ2yduPq1x8jfNc5H2K7VPrAfvm5Z
dIFAnztTYnio1TCB2DpJaee8Xf3VR8cIZOmxMt15Y6D2BC8yt0CIy43FkFbjfPQlVJcIFMrZspgQ
d7NSgLrADeWvN8aJ3U0e9QcOGOXgjVocy8dL/lCYaMWvovf+Pi1UsUwIRQ7TWcy1LH97+ARZTj94
sRVpseWIlNJWPjXBf8UvjCY8tVM0CV37EPev4YOZyt66UXWnNCNwQo/ns+N90qnQFrn1TS52Mq+A
Fhb42uNqIqwmx/TuVEJr5USBCDvWNvkoOZ0ihUl4RWtUC8qvcWfHaeLN/NytoyUZ6xvF6VDRwUL1
TsLpQ6IYnkVfWUeuQY62FiSQjX9HJAUh/RO8Sh6EkErjjlK/Mav/cJgUYsPWDlwBAIc9pK7iOo7q
79OH/gTWE4p/o+4cRpcgZN7fKE2/2AAWc7B9jLKJf6MtVoWPL+/pBRbPQMYGor/7A4kflU47FX0q
tPPCsQpR4vLHCYkXeIGm3+FD84VT24ECtFGyDmr5zs0FlicJqos7zIz+BtrPXdFGGfNcdh+2OHmy
aOXjFw420vW/HR3haC2ghoMppO9w9js0iNbyCv5mLbBWhGDcf5cK8KZ0ovOlwBdKBAZK20lYrLuL
IkdpVvRd/BtsbSZ2H5rM4DnzPAQXlpBr7qB9MM9xw36AY2Mhs+SWv4wD8R4MplhdGhCraZQq/1oO
11P/KJ52mdg8+WBC+hFx4+zK757q+fOu+Zl95fuJlK+5SRK2i4q86b8/O1PlaNxxTkPUT/yNUF+x
6PFo1lLRehTKXLnyxMUVPP0TR1kYR7557oKU1ikp3OwtHZ5vHbAhLRKh2tutphhejNpBrxLCVADI
vYTa2fA1Ca15SRVwktwlMUv04kI3c+CcSkXntt+C6G2aa9bec5UxAH9A91Ns9zffrb6lrdbnmcJX
76OzORZGGdD589K0/vwJo9wffzXcorK+jp/ALZJTqsnMVY2qa4NmQp4CHJIZ1wBvk9nKG97BR+Wz
BP9dniFLWk645e9wyEjdR8/ZfHVqAEpHyWS9N9OKD5Uhcld6+eor+UEeE76zVJuNh4+32ETuiH6S
ybfV8WVoKP6ncIRlZXlWa2sx2efJzTjae/CqJPSaH9/EkzX6Jth8ialPgU8r171Dzzy6Ka75kmOf
c8EZJaJSK3SZA/YajxRrl7fyxF9gCMJiWmde85vtGpnDawNX+QLzmKcYAHy7OlEVX4F4xmrmy1r0
VjX+WlAu4G2bEg5yZ1/e833fHbfRwOK7wNylT8NrfHX42kSwVsAFL5VwjHGhxuTZ2RHhDT/N6h2I
jyXFFo4qU3DYVBwHnBA/+PmqZpxuqKBrExb8uZaQ+z/X+VGSM/8t6w8ZM9tC70q0IMWO2KCmSrE6
2TP8ij5ejm7zgtq6Uzr2HdmPOES2rhgpf2r7m97Jf4zVM10Om75sYo9by4VVB4NJ/oKDFX//dR8g
uYBz+fhC6YKhchfbeJTwCjh6uaRAaJEItviuod3BYEvcgxPbiSE5csnmwXEF8WLhsgBn4GNbc6dE
p/cR7eS5DRf0T9H0b0EbD30eD8x6DqViFmm6IsUV+JH21scU/AiF5tl0PlUtXw3Op7z4XVzDJLJf
CHt1VDwjqrGK3xYkRodTiQIztyhVGvZA9zv8vhibACmIe/ES8f56NSGBI8FpKj3U+Ksgplc+ZvKm
CzpjzLumlj5zpSCkIa98RDRIwHUecSURa/JdTRmvIOJ9U0y3VfpPDvKfJhEyi0tskpSOjI2LLxVW
vRRgBcOfz4CboyHOV+wljXuKHcQ2r4OgZe4Gm2Aw3vHLZw/Efj2wsjnFKdE8zJEsZr2sjhi/qDjI
AORq6HyDDEgTzAQGKhkt9k9lSSnpZxCCDkRBonU2nISEm4qLI/YdAKr3St6vBKz/iaVVHYym2NdX
9Zm4xbjYVSKgxXqM1xpPFkIoDR138UHu2sYvngOa+Qzzega1I+Lh3KOWqsyh3KrX2i90VkZBB+1j
8df95tZSLdSSYGfKnIFzF8r5vmwAvBbyfm9XHUjFtYJ4vpZV4fC1clMTu8W7CoKXEXTOmyTt9oMc
IjggnAZ1+T/bpKgR1h0y42mFwkduUbAJct96dL9MMF3rnS83pqZrQcDZmHJqxKWXJwcrHloJx+Ey
4gzbt36tLH3lpvFhyxEmMTny8TKPllNCwMFgp8FDMRRfI7l4dsevATl/Td+nbcBVg6y5wI+fOryr
qfxXYxd4PkTyQtxn7XbwNQ7sd/PA6Nbo3+6WJPthwEKWPaOK0IqtO0cqdyC3zTdboF/MfisFlmDZ
BUwZG1LWjFI2ZxmuBkpT7tYHnR6zWMVmtqKrwrQwA6RIReEdPDtCu5MR6tyysHRdUIWjBiJsQ+0k
Sur1d5X+S7YR3mQVd01xFmPF0Q/HH3fvJ6U3yQin1jFRriSYZNSTBAThuZ+0O+FSSci+1LXLaknQ
JcArOOF6oxoj8TPpS4LPeECiBOPwI9N3DaZVY7W86PFZCHY3Gz+yT46STLvIp24N0Jcbm+K0DxI0
RrCOENrEiSMnN+HRpc0yQVPP+njnAVAyWUwnncmH/0ZkVe9q6ertj3F9z6kmtt92XHwhtxuhNni9
Dzuq6BfrCS+xiGZNN7pcs22YIHIDYVyyeEo7GsuxgPIDGKUf/wUkMO7qhjmN3fHGICefw0zGQ60X
MLzZXXKpfvcfQTWWd5RthxKeI4fnPFKS/B6RuqLRM6U6z8qTJ4yQoEwQY+oLdupYBXYaXCNdc3Lg
I3XcFblt4zqRggPR9MuQPiorwsLpndlVUwpgWdDTjQy7U9nG5zuIiCA9yYq37ocTN8arJYr7/7w5
CXZuDt/O/eNERaPAlvmrSFVa+BIEjmrWy6HGCOJyVyBFVNp5CZ009IO+ocWNKLPnMTx9E/jo7IoD
1DcHrojawaSE8IAcdWkVIZYRAaSHdRZw3ZASYobwuFTfinTmN+XS69eGDhQ8IUBECCGrIEBCucvm
eK+rI6m+jiypBxFaLvGpxksGNeLV9uxPkpsGReqpjZ/F5YpZLpW1I5YC+MJ3xTy6xADjBUkpILVs
ZMC9DsRkA2D7YQ6HR1as+qfQKurPWEKEdOh1AMo081Ye4ZETUsKE3W5qCbwuV8jvTRYFAdZCZ7bV
s9H1f+Co0F1HFvb+DAKzjz5aLJFQKmzh8BtUVT+XisfBD7Bz5PblAVYjQD4zqwaE9FlRzjKj5Kl1
QiPQfs59Sv/qT8cZgBeRc9wj8uYcg5ja7k1OrOURoevnjo9e9wc972fQZVKZua9Tn5ufGlOEa2fu
SuJn1ZwxiUE4vs87rkcZs3n6XI+Kv4jp2iztwpfnGAPQUbwWMUXtcCD7N/WGByrav9/MgeIZ5Wle
m6cUvNcqcL+JmV4KSilXMeCCv/yeFf5MBsfacYcRYOpbBM70KOVoDLZFvZ8XwfTKdLB6GKsTXYcF
2BZZ3LlVddTPu2rn5lv+X10XBZQC/DTxHOaYRAPbaU2W0fIajsI+bagOEerFM8k9zdCw/lkkGhYw
uLbon16KYFDFUp0qyRRie6nKE1vQtcXrGlaRjbXohYL5XxRz/BRJSqBFe5ACv5rjOKLPAUyfdCve
v/mcyrUlhwNf0tC5D8O8pS9RBmOtX9WUkISlYnG1DEQVpYvpIIP/CehvxNz3VyKI67uYTSgWjTaY
dxZ2Mp6EyNXAQQ7bInb9FT/2yByR6jBQkCPkWvwrvDbquKBEAXLZf9zVH0bKZV7y9T06EcNddgMF
NRfAiQeWwf1qe00tIZiF4URYYa7BFUycXlxVoB87Rjr379MhNADrZuvB8NmUbA2nxHN82Uitgkit
IO9GzKJ2fRBuXzXec/rFLzE8QYqLMWAPacAJJ54r8GHCPyi5VtnAI/lVxlR0/sywTTkyT2XMF+md
J8OHg0C20g4rczjsrLu8GuJB4r4jhpMU8kSpo3Da3Q7jwzyAisxGfewKAg/gCyGMO/telKfvHGHe
R65Lt/1xK/PY57AQn45Bqe26SxjYdNVQxmcd08Bt/eJwjKK3xHZFgP/2ztK+ZfcPFDXIIoZR+Su5
TDPzXmtUTxqt0doLskoE7B4F2OzEFaREnXnNXqGv5hLoSCzD2c+MrZGq6S4oW+ST1NS1FZ0aauVA
Lqdk+1fWhGZGBVGJheEQrkaav8Aa/xFk6fcqlNLhNcufPkmmIvXEBfPkS4nCWzoTr/5e8CFnyEuV
dyrvii4OiIAuShCxIf3A02X2t2YUEcfHPjK3DIA0ZDcwFlv8u2D3Atc8obD2yDfOIimovnR328Df
C+fdMh/iaGQbr9m5dc6/cLaBcKnSlUZYbgGSj93/S2CeBNRzkcitoTM7co/LENFhtJSBwqlBOwm1
nYIRG0wK7Ct+4nAeMcV1cfNypubzRjLYeelGPxFU/uJ7Y26km96SdqmCw16J9GaTWiCfUcSPBGrk
tY9ZsxFgggTbaOaNE+lKxMND9Kg0npSwBXjEpXGlz+7f89QXV0cSYSiJoBoPKSKTd8Wt5STKf9WB
07qKttGqLK6wY8w5e2I3130pukF7q9RDEG7G2YeV1YEaYLpnvMuPiWigVhWxdCgf7rwtK87jGpFf
g11p9K7QSKTSKvwB8E/iEiGDd2YdyofjT/s2GPf4piAUNvqOh34OquPRUzQShVOw5e1bsxAzFGGY
sTY46q6Y+CSIy4kZoxLTpNKa3HW+5NLxBV9O7MygbjQko1VIJCnmOQCCpzGJltZRirso+55lKr2W
An8Ms028On9c1jyMelyNJlwrg3rqkS/0VatsioP7JEOWbG4rCupPaq58dqop+JSWzAyMpMkZShQy
3/nmN0q9aJsO1pLuUsnaIYzp9CjP6PFynrfboTqMoMThrxXz6ko3RfWeYUa8xcgirs3SyI/07mBX
d0KCEsF9hE505cOGGiQ19A1CLDJvNYx5M4Ox1yssBG+Rz9giXumr1iUgaxtrMax2AtgCC9Ltq8UQ
aWrZ07kNvyBai/PTj0/0NNEiGZ4EgYKI0DGEhEfCx2vV5fdwisz9dxL97+yDduu9ruk0I+KF77nY
QJTZYIgRZMiFvn3+GVdfqxzkzdihX72jbXRgWerqoLsg0kMfhMbxh6tWpXzO3w2QMzQB1I1dIgqq
vU4GKUHLSOHSRdUsBuCHZ7AEikRHIJKVmqUqH7Sg/EM3+jYNHLMwAK6m9KL5SSTFc96dRPOWkNDI
obb7Jmm5ERBQPNmfzWHJMzt98xlekGyRpNwSyFxuRX90Kxu+TvUT2fifF1K05PzTlGrB6DTvnk09
xexA232iXUSIwyG9wqf16umZFg5anS6vQ/2dhxynAT3BPA2ErcysBjwy+1Aj4NMbqJkKQY+Qf+C2
kfFsrgzGryDOS6iWxO614boOvgc3cmECEXif1Etf1hJsFQiT9DCPZrWyfAv6ispsCCmvPITIUoWU
Ntq6vykRI3aTIOYLVJby6ORsz1SmRNPUHL4VPPwKbroQJIC++21d6Jtx+694zFEGJXoFm8JQ7C6g
jlFPGvS4N/tBSrFNSmfdAm3TRJxDmX+Fq/BIK/S9BMeQLMPrgzGU04MC6em1iHh+Btf2LSnOZPt/
1VDzRFwAychdAJWJmmpo29Ba3P96EzcufCzJW8mjtI6wPfW7MSNRcCZZHu0dXKCMQFGfLXHZyIzW
GAAHm9powbyQvmzAc0pU1shpFeM3/MXG7pn3XfvlDqP2AyZ+ICmFAM0G1Zx41ahbaBaTSF7PRPrS
EEQkb5XFMzeWzveU9ujKdn+SXM0BSw+9UWfzJy+eCivKIpcUWumjmbKENgr2biXRtxnQ5KFlG4rq
wGbLCRUS3S74N3I9qI0d3AXqrW/jVVz0oufg2Rb/EGGoXbOqZvyzT2sO8QOynGS6HzXJC0FGlGAF
EmWhGJ/y5EA8NZELiXGutqh2ceghoIsBEo8e2r7Qfr6s9J5SyWPxB5bMZADyEZhj454IhmShjXVb
UzqzjkX6bVPoT1xiYPAE9kCfg8gKqyc/UxKzbHWT7hVp7eiUm3j+W8i7NavZoAB3TCihgLYnb4PP
giVwjjvCJD+rSNLRm5OlpYRa19XtAsy7CAVLi9/sCKBkVxnaTmpqVOQXVh/pRHgf01Pt/orUljcF
C6dRASKLyf5tLCA+QSPWGxMqbRCHf+WfOB5oURxSG+AGYPO+bflGdaq9yimrUjRQEOY8NY7NCqF+
UF1MbHaeY0HOwzJLgb1l3TTke3vkvnaIQ6WrQJQydeJmcjlgf8B26+r1rkUAP5gBezdQNcUDsNNV
CZpO2eWSdQurLdHRhI+YpxVCDT9k+/cjEAsmC+J+DUaiUnp+215g7UPg4ZQi36fx6EtGU1tRpVnG
T2XT+UGE1/ag+2ke6jrlb52uY/Nwui7fQ+85ue3XBu4Ganb8vTK1uliJNL90HjdyrxCD4/aoqCc+
jAx2cn6a4LOO50CR8kN6zQsATJz2ryhJr6ekmlf53HjoOa+8RsfgcEuYh4bOI5vGJRwA8Z8LcFKW
0N+9H5y1/0uLmXo4VCpwlTAswi58Zn1USgRca+R3g3YNxdX0W9aHiPgQvLK5zsmW9DsjcZ+RXWH8
2Cdj4fZWNLYb5XLaoAolcipukk308Ju7DQgynM4GEaianUD+Ty1J0uxeTscUF5E2a+oq23ndsU6i
c6CM//93WLuLhw8XL9vwalmOlgNuN7bqkXj1auIncVp1lOQgewblO1W7Txzn3W018XIpvlHqv7Ww
a3ve5YJm2pS70fR10kBIhbK6mvwRc6dN920MEgKXXJTb7YWdrnPmqEZ3dk0UJxpI+O/VlP8bqZxz
TFOJPH1cXwL8rzvo8ujShQEyVG6U5Q/3jGU551CekwdO5uM1p5xW0RHKClEUQApVUzporq6sKvig
jfdLvqwcdXFrtcXYsy+3ADh6gB7FCGmI+3SkNKp2E33WXt7KSc86Q8juTYipDc3TPYHu3mNeTHua
X1Edrsf+7JZhrlTfSSrDl9OOC2nCwz9fyex1pY1Ku6OXOwyX9j4Ye1veeGzk+x4EDZOPXvds6bwh
zCendP9lTRoBbLidxXFWCkUoaPXvdVVBVUY/POXE/5S8ZzYIwlxyz0px5ysSyhdvamRyai9Q92FM
1SWFQtDijMVE7uZNg9RsgZJLknIiGCYgZO2Et5nCCcC8ZNmGTwhk2xz7m+hmAlHWDbLgkIn4KNPR
WlulYZoeU4ncwjxLXx691wAIRsYWLrAXqxQgnUqcW9uIxBIs5tVu5oMp4LTmJPRYm6vcOvba3xD1
MY6eJc/Lg1ISXHt9Wbv9LMCvY337tBuLuG/WQxA9A/mfvGs9UeI25sz+NkLrtuNc6csW6ts++5UP
nX9WC7E9NDpw5d0G1HZ4q0pF9jo/6aysPjlxi2fh3zNdE22cgDCrKg41MbEPHwHKTXwMYa1yEQrI
BF2v7yX82nggR3PILGXBMhoyRIh3YQjFF/8BRPr5H/FkL3fyzLVxaugDiXfkx9ub2AF6U9BuDnRI
ABZgvqFdx9KqYYbpl9TlgNlarwmkW/gSJ5ziSXRnrF1gBND6OntmkNRgBvslW4o9jf0ymEW2CIbt
5G+I52AJAJpse2Q8Vure2IualKt77jbAfZKU9Q4z58oYXVij+NQ9CqT70TXxe2a6CgGmhxgAmgzH
TRaHmS6MmGupoFUshA6nTzae1EG3Y4+YZLca6IVvCZTOEoTPoxScGDwN1JdLUgG2u7/BseCAyqyT
p6spXhjivJ+6SlbZkE0yj7mAOl7pRlr/mPiGZCqF+G7dsu3dqRUjuU/CVazDWt7T5hARDJMpUbJc
KUnn6uLpwNZ4Mgxeafigep7JWQw+lTZxPknZRDH1c8IcXQ0s2Jo1my/Y7C4xFmtVlEXfWPonlkIC
RER1oohOKJjCQBaeg3nhUByRg9vIUBKh3HuX+75am8YgeMrbUuT8QADRZ+fakNGSVqfrEpRL2kLz
KWFWJMBAIeNZiazWzNeK2Gsa29ifDu2ufpGEUQp524mBD9OmhzmXNiYRpySGQPtklH5W7/11wGc3
FbnPYSufTvTZDJpW1Evaw6H1uM1Bwh4JazjuPfcA7toprjZtUJel7hFcdg8GeGy6u8MN2xpd8SrU
nTUkBi/d69ij806VMppA9xe0J5HHFX1+0bzHAr8Dofiaz7b5j3k8xa4RMHgx4iEjMa2yqo1iP1/D
xb30sogp8A2yuWJL1d0pIeWqbVA0U+kutsOlmPNYKBcv7cmO1PAZrOtZMyubV5LPKeBedEzJpNLz
6jfGlxAppymBB+WkYZomoFqeaY2OFELc/WEsXHfIZhK12WqT9Jl3dwrqkGX4s9rrVn1Bv7pcEyhU
pzWq5BrYYnW052W+fLmrXeHwZcXqlsQU3tRkPSKY1IheW6+1PNEal53ZruJqOwbagShHtvqDcwuo
W5fFCROKJrObKhtnQLxALNFlsKd2XjCYwxSVRsR4dkPlv4p616JQXI+53HPpe7IiagFdfXUAmdrx
28s4wPue5rsIrzDr6AM2zfiG7q3/Igjx0KkA/p1fKEBGHU+vbAkhvedc7CJf7lAGdf/631kxVe0I
hR78fFja2JjhX0ICxNodrBOQo5IT/n/ngCIdgPRir9QKkIHZ1AIxotu+NX2hgP14M8hl6VIh3SMC
NfEvTTMX05uVDPLB9mRV4CmMDkLy91jOmcB/AblicCtmg+L/8FBYDaSv//p8xNr7mmaj+r9H6P1T
sy3mJ3thavG5bl+6e3g8XMLwF/N18ZK62Rzm6VLWy6PHzQSTzu8VmYjVdtmfcvScfrd1qaEuwAOz
NVtGHUDbagheCQQhewKvsYn6dZWfMkxtXH6rP3YXZlxPWAI9Go7Kp4ryP5sLtAdh/sb2NNRZv2nN
xJtReic4pwS8wLmS87yfy+Zd13/QC1RmKkPiiPdHQgax+ecfRiZ6rd7wjex9t2Cv6QgNMtnVwYR8
bK8VX197YwMcIpcuHkcN7ehUSHmiXhxT+WWC2hWxhZqD3TTyhBL7nPn4di/jvmzpYCLZgRMbItzg
SwBXQCI4+F4HuqiBD52G4XO2jc5s4fFazrlesUdkaqd0PcAZvP/F9Rxpl5z6VBQllkrOYjZJMrtC
YwVakBhF1vavXb2XXoYgYrocM85EjP5hrQ6Qx5ixdbH9cSWvdOj+DMNri45/3NHmcWoOlyql1aYG
1pJF2SXLUwWq1wrUITEWP9sGxW1dmOi61a76PXP5RzLm8/KcFf0WZGp9TNhJPYupSpGghkkXbqvy
MAPw0kB9WF160gzKZmDr2EcmFfV+krUtgB00G6FdLVYV29W6SUWJpZ5oB62fwCzc1urb6pc0j/6F
nqqWEmuk4jP3534S2NgKyasFsTXVE8/z7gFrN9xCydNGNeBhJ8l25SCG7atc5zLOmu8R+X0ngWVQ
x+dq+bOadZ++iIZAEFF6ruy3VLy869PHuXmyylp0DJ22JOrYejmEj1KPyEJsilm2E+bliDpcpN/A
GBfqOCpoBMBgJgFpZnmWHcc2iMJHSawI1CpaxUO7iN9LAE5r2zXn2i0+1RnsmZFiOdzT+9xtxhZR
Y4hxvDZu9VEDh1hlMyV1kdF+0Ct5ipLLQhhXdhQ1G9F7RlGo1NTRYeBPmoUYcwc7nR3h4a2oE0yX
jx6BEoab1yKxBL+wWGigfQMJfdV0eZCrXzqhJJMaJl6S4cFfbKyZW9GjEF/iLZvVc4MAHV+bm7RT
y+csPx2Rx43F+ffiDYuI4CpbQsoAMCpMoOYHbWfLepv7kdrBrWa956JAAEZH6CWoTXL6GxMOXd1E
So+werAjRlmz/FjzWtANtBh1Lg4Wkm3+bWhVw2pjQe1DRvhLqbEWbdnfyYKmXYT8Tlyma8eyJ9E0
HI2qrNsqj0EOhc/ytSZ2Ad8lUHN0N4Rg4sXdQ8dZBAnPV7os1Ri/kxnEA5mVI5LCKL5QsGm1CDk3
1qaOnxQ7sCyKzrKpqeGv1S6C5CxRlnv7rrvN42M/CjgqeJtYabHc0vgDYV7NL/kE6q0Wt2Xw6vx1
2wFtmy/pw1qfhR0wHLTo7PkA2DdhpzJ8vaeb6tNKrtOVYxfYl9Yah9I+CLXH5zPkCgT4EoUh20ey
3p5TgRlcDACczZGCFJvCl3Z/8cKEIMvnOnGJ3l9SfLlNMTv4kwR3usIJANe+90Ct9hzlWxLs5E8p
3WTVoXsgC3GS00CBPuCRIYwvulFrr02bxyB7sPRMCeMe+aQJEcBrod8cg/82E0J23cpHXhJpg6ly
xVDGLUOJFm5v7RkdQVvAks6WguJy+Mhlq6EPky0CzajSbROXW1nx8hVIicr3ZehZLYweYTCu7S4d
1kMrPazpEH0iYV37STFyCEFz6rjzsNzEBT0Sg/cPdrI9DS3jhwYretBiGlv/fR0aM8bXJJbpGA4I
89VORl8lpPc4GiNP9kXh8pcxw39B3bIP3XNfibQRcjEla+xa1aRYRwuYTZeZLo4bUE9O4fLmKuH1
FkGeXGAOd+0oA/Zd3SUYvAf6DKOKWasQeztOzu3Vcc6QA3Iadd/IHwMITPF742f2B3L5MFgyGrlN
nBQeWDkDuRyAGkLX2K5mACh4M9Rba51bA6R3DcqJGGl3wcW3Ml91LScXvqNWM2DmxLjfiMXReY2M
/MMRPcb3kXEWF1NGW7GlSGz6qCfm0srqFNEAZgcUjkqQ6kIuLIoPXUAa0mZonHY42TJNA2V0KIYi
/NoGCYri8ge+bwtfkERBj/KwuzvCcOJGik4K2h1iXgTZaoU2M94+m4UAxR5eOcFRwvKVys5+SeHc
AmZY6AHI/ovsh1wp3kmLgJHA5WME3YyviFhrRnlpCl2BmOjAN3emVDDCx6QIHUyATV+mdm7wv8uv
2L4AIIzPr8ThcejakgTLq4YCT5R4fEKpPQJfZSiKhUKguGRHgijLseluZhMO8svaFSvbRaXs8onJ
5gg+Xu10iaPDEMkk5DatDQ9fMep7HyqrqdSk5hvIY7R+q0r/NsQvG9TQR/06+7RCSuIHWmU0eZZM
GQCKvi4dBGTETKQGf5bfvGMcScZaLw3eWTngmNcLwpsSvabp4et8+b2Pz4kNQvUCN4LG+xcQKk9q
EsONf01HfpV9pXMWOK+SwiAfh9H7ZyPk0rT3TnP4qPALjCvkJGd+G3MSZ/sZdha4QSugDX/RdURQ
+uI+3OIJsRK1EjEns1W2PYhh809n8lja+TAeltbSeOwTFqr3wB4Ydxp1i6z+8NRJr0a4cZsWYIdT
6u8JfpX9B9bkz1TG62pPMYhthOejAB1SHNpUsGhjf80Z7FGcSJL5I1EjfbrCNp2VXQWv85jBZmLQ
qLAUPPOEqf0NAPangQmUBVDMOMDdSCZ/84IEe3iGnnWK4Tu4iBvweIHGterbEWTz5r9nODhtpHF0
On86UTainUU3J95qsGsQ0GQmoe5e1IL1YhhVME27zR7qHdZs2drszYxLtWX3ZNoqW//GFrmDW5SV
tHBzaHA4QOv26UBek/RTHaFnzbBpUbpcxKDr6R0C4Vw37UILa0QUyZTCLwR7biTMFLbu/+CgWKEC
KJr+jow4w3dWPzp/8Lmhp5otQSVTv73JuRwRVztmQ0xElL5zzm/3MbokJsXHAnC+CJ2iwX0/onsa
Fts+3lu0X5jSWIvvzv7+eopm23729QX9N5ma+RORimidkggelHamHBd9wgkFUEYzsGrS7e6nN7fn
Sy5zpRWeYtZ6B5b2PajAoEnHI1kCjszgIbd7unnAkXO8E9D9mvwRqFOj4gPYrHGV7rb6WgfsCCm9
VWX6nfGxzFY1MNlJ6iAhCKyOhcbzQv4wRhyI3MeQZRH30HS6wkK3DWL6K2nBpzr2pQWuWODabofN
Oih2F2xgYlhTgIcTaBjBR0FaWeWl7iraCYW34ZlP6SGRNsPeHhuYtXTozZEErYUfZr0jkUOcReSz
dupRf9IKwZa3hIUv3Fb/ZQVUQhRr8ABub+YuQ746luyphuJrb3wsYPiqovZ46UuOFJRfF07eX211
hhcAfudRl3fLgnVQHzwsO/6HGtJyw8eFFDzdz2xJyVt1ZOyLCaQ05m/P93UxR/cBQl06bj4dWvfV
2yC1OH0Yy3FW516Om/hDD5z1KEJRzkpjj/KUm3Zmd7BcCzHZzFu4+gUD3iqsFHs3fr2f8dK52gWb
GrXq8Xl1Z84VpQbtSQy9fQftyqW5PHwr6jwSHG/tlLY4WNhXnGM2F8s2WTEHQJ85WYtgyt5Sbe/8
o3QfBcPgeYRQGeM9sBn257Fu421GhK3OoysaQKP6s/2imr3ASjI5uoYAntvKVZnHU5o1tRkGvhR0
XcSplx1HNI2FGBOkSWJDiyjLSn1CBKi9XKvyrjoVFu5bO6FT3pzUSjcrKHOpyR8waykM3tvqmz/a
o0r60JPHW00aJpjaBud7JJHswSqiy71lp11uW28tlCip7GR4yd8whHXhQonjNYJyQn+jwP2QVTbN
KQ3qKatnmOvH1+9xJQ17nOvsrAvzW2jlTzHHCu6OX/FNzJYz7ArPHOdaOJcsD1Ky8ZJF9okZzHk6
g8eDohjkJAKCXBXy0lg2lfsAmMoRP8MHZglfQ+6GGg20i4wPjSxOsnWdPt5dKqPxxgzeAepDHZP5
kC1JquEeRNkZeeZbaGPwdl4TSjjGPkqfsuEr3NrZgDE/LmzHNE14iwfSs+911vxsDT5i+29F0Gje
NAd9qAtJslUs6OXokDmu3wpERujzFByohIl4NPaUj2rWuJH17oxHV7Gw27sT1iWokkW2bQhrrKXN
9cb/l3c3K2JNERO/pNmvREbQznVqFP77pGDfrf7SESPBKFerpryAfCPc51Hicc/XE2a4zXj7eD08
yj1/Sp1l+Cnjof0WTbpaYKiHHH5BacQYNyb3MezboH2XfvoW2oc0PfvyytLCz4FGdUqJLrWuyGT8
EAok99gZuQrOWBkpP42zSTYo1kMQoRGSmuHA8yqtW6b6HEugpZGveqyxldrDrwIWiL4XMvGzHptA
1FHaNhZGpOww0Uu4j59XjTlKiFH/McO8a2sKZrQXEUAM2cEl4S3D5FyO66jmR/cHhpfvbme3WDNH
iQBiOLIq4hM9e2tetgM7/fQVSzdV25kWRK1t0D08ZkfhZyzNR6CMyi+JJeEtjJePz7CTpRIJMrfs
PcZ627aMcO2ppJiyV2BAr6tOKWH7aAzZQ1nAe90qTYFG/3VE2WxlOTEFtrhG2ShBdvYhzp+acyrT
oNkMsbUyCkQPNXT5o5I5h6CjqIS4ip/qcPrOrSMLD+2b16bf0azT+pSzr5gyecE5r3H0UmSv8dem
RbidhYUR8Cx3buCWytCuAIBOwovlidNlRL98kNxTh98F6fv5jAtbdDmpC/SABTC/O3Lt7A/W8lqB
inRHbXQZ7HypfSypvjP/74EJ3sne7eHrUOlvOdIl5le/Dj+RnDFmwTkC8BPcOuPEHw146zer2Hli
YHtH+3NFNRlvIYICU1bQcTRyZyX/sd2Wu2CmM88VMca96p4tpRWw82ui2j6U1+p99QW/1VMlwIyy
WA0LYiVtOxjkStBf2OWuBoyT65raxl0KvQqhPgYc1G4WJKdLvVghixWGRUY2MeD8oq+vTuezYSdT
XgE5breTmsewwSwzTrNF3Nshu0ekD+3nDDSZ9woxXNc4MqiXeRwlw79qWp1YPiZhNWlLF5evUaeV
xCmt0XJhPib96szGvz5upehPmGzSslE5657GT1SR0q7W4DPAkI43X0mk7KarHagMn4w397oP+Rwh
9XnecGLvjBvw9UZeq3OkckANTUnR1vSd8cbNx57SVEk6qVo9qoL4W/BjcV8sQyRhr83Fcpr7BzJQ
+1lDmvJ10sTkyriD0ryej2QDBi/w/erU2pOO7WKkucgCKbZZfaxiX3STCf2yPe64lMWflZGbqyZH
nlahQ1eC/mZmZYl5ZIOv+2nMxT7td0aQNLE6BrHkhK7cHgSJ1jkEoa/XcUFNa6NiIFnJYLjTMyyN
IiKRSef+YX4FWXRa3OXxHOIT64Tzm+giUFnjRkUnNO+xerPuu6/YZvE3sQyDxgnJLdQYIojOosxu
GOUuFg0+PMNJQ9Jd4KPjSPSb+wZTsqIfb9Xwp/3z7vB+hCmXWX0wlmNjwAt8AOxcZ9Y0REO1B54B
379dZ2TO14QbN8hKddKdEzJ1GyUvVn0HBqKNG8/WEIP0dNlHG+7omSpJy/JauB65iDcCm9ps1mlO
E5RdH2g/GimJVusw/NOOjw4TVRNm2vXL6X/ISnsERLRmbycSC/a1ULGeEH7x288m0TrmI/9qpbYS
wwMEww6WuPjGoKHV0JOnVeOe83+/f/K8p39sR9CEB0H7nGIe/diKixIYchnERt/AGD1KpdgGrr7P
SV3esKG3Zl/CRyUS0ZIJ/yh4BO0AGJLmX/xnka/uK+KFUaeR6lW+DYn2gRkAubT3yvUzlbFVep4l
ogrlXAuyLxBRXMhIGlTiz7Ic42KnUHRxfy8eUYRVGJJYhLdroImVHJe2vfmI/+8KOmxt2PiCzFxf
qREswUFnqqyhuZyEJSpbWv3T2YZ6zhTORjVAbx2nAgYrbuYKiHCo9U303cjFtyQGUhoYvtxdBJd8
kSVCDg1RriQajIq3Bd4XXYV7CkcplohLEUSAWUe5PNkveORGAayjWmFs/KdX3BoJEA+BDM6Xdstx
+v/oSP+JyF83Oz7HlJixk44rSWEGPyRbGqa+ZONXkZIAX4+HvxKdTbfU1CFweIwl/s3QFsgUkFWn
QQJUMEabghZAisVbtrqo0nLM2gtFiumMQ3svkMR7tMD1B2YZ4Hn6LDukQMfWHI31d4rG/SfqRVQx
AwEi4NBmFrnouKjnc80a+7tkVD1NSu3KoS/5h7BAo0Y+RjrAxX+3o5m1i7WFSYYpg1I9JBICH8aT
d0vV+xVtSMwTnj27Mb8vMlydwPNu8lD5tU6SeT304GXnCgCQNJNn/hVs9TCzCk6wdspm3r7wqdAo
S2NIIMWvSQHcsOaE6lJRTiS+7CTkoaR3cUgvHYo2ftIeSQ04NeocoKpuerPYReRz6tL9nQUH0LKX
/++uXLihGXY1dwP/Hfb6h6aYsQ6s2G1Bz2dgFWX9FUEUNaxOkf/WMaf8EolkAhsnGaDGyk7aRDEF
uvWOtY0bLvemBZnuOq3H8/jicG8Q6SwBf3408tgT0GFyjYGC2xmn7LpjjCt2Zt0tzSI75z2friUs
I7s5wGRa8jHiBIQK5y5u0SUClRKGNdG5neuI0Td/5zkKDE0i7xR+AiVaf8wVY246Wic0BrMb95cI
hlY54e/qSF8Y8SwjDH9q8hAJDFW5SEXzFV+Jozhsy+8IMg/XfFgznPEN5K6nmjHTfOfIOVcJfokX
6UC+KF6aDrhTfQpOqGXJkZsFVEk4H22wvnn8QPa/wIw8JJmrCjPj6b1F32nMb5JzrHM42ibgrSD1
Ad+/zbQD8S2R12rKoUpeIkxuGCeELS6xAVVkCi3kRgKoPs6wcAELpsGuGKrJis0PvrBEVDD4SkpS
OJv1z3M7GTEx4+RfIy0AISDa+WoPcgcRtcWfXhfwbrblPc3aYiWpdzfQKiRjVS6HE+OFoPI5YDKu
tfr2X8UHID0PfqjrA4mvMHIsp5u5+Frk74wyTvX6vpS3VvEC8haVkplPaw5eoTo+IjVHqdQPjZmJ
u+pTlYwRzA5QSNea+7oFcsSMFAlQpO6gAIWUuaMmvuG+tucDlFL1nAnQsUm34rBeUXS6M8Lq/bWN
EHVe9vMz0zcjeDWbCd+lKdF3F4vjAPLS/tsy/omgQgDYm+2/4p1Y1nJi0RRJ2Xl6h4HTisCDWebv
hZCPm8AhslqiNFtAmi/bDitO2F04VLqNoWO4UIWZimJ9uw0rMudHNrIWCT6KyHmcKvED0RVuFuV0
DK93qBA15pIuTCZFjTWFlP6k/LS3PP24jIcJVvRn6y0p95YOEdi0HI7jXzWifpl0e9/NcTEk+Koj
8FJLLEzebkKA5wOH4sMmKR6S1kC6WW6j+CG7+Gl7+Xgbj0z8PXr5uRq9RR5QlgvSx2oH1I6sKQ4l
gXWftUzNYLHrP8LWXRXfZP+MSWOpAjoney5tWfg6sfYXPJ5koRD7MmnJPuJ1WH1A2J8/mc8UlJQb
cpL9cwZRPAbjoD0ZcT8pIcJQLDtZIWcBoqJwCvPDVkk+ELVXpfBAGKH4qK9H1uf9yZXJBmaSakjf
PELfwzRkHmrjUsc7yn6IpvwNa0+2zqk2yD4rQtDntsn6PgVkNCCOSICUPDfQKIWcbMrQhTNaoBZd
ug9HKKrtvL8KxFL2uwb5X/JevurNT6ncWMJjz8t2Uf2fpYC6RM2UZCFIuXoGB3zTVC7nmRKvDDj/
1n+/Yqsg5YJ7IT30J4l4jm6WqRlOuYtenP57TYz/z8VC/IqQ0U7B1rRKyWRqI6PdGOyd/H9TIA03
YJehvt+TD5I1DVTi7c4v//VL7AXz1BQ088gr1zsf86Sclvb0dbVI/Z021XoCQA+TMfe0M/nEVTTa
m+73PS3WJ9+KPx1nRuKwTVH/dj6LrECxPtFA9w4sIu4QyhdrPSToG37ep1d9ukdP8LbCoD81FU0P
MX1XAYm68izqhdjxo74DjQFem4RRbGiAQ+dnxV2V2Q5XRlS6+iaPSRF+X9SYD4k95A6BHd92Z0bs
G9FjLwWLPSpcBeJ3L/EY6/e8tVHvwkAkjwg8ctqzhYEktmK1RM9rCwW/2wzPCxqMXaTk+dL6jIbZ
mPTgCcYezgaAqd7rAAIq51NczmfRA426VvwUBNVm0ojRDNi/Z1JPfdEw35oUqrjHMtp22zO0wAUQ
bVaJanNB2VfcIWewEEG9ihI/X2eouR18ugn2zTqnrpAj0+mS33kG7cq102iuCBN/6mOxseAsmUEq
aIU3CCa0F4+bJLEoUFDghTtJJHCed4KXknDacKSorWzZb2DE8YeSV4U7aaRm6i2quxKEL/I8CP3l
D4gFNWyW2kFAN6mTXSfcsEiOXk+L+opJgxI06unnTQ7m2CEOGjB6gQ27qX1WeEBqXm7xYhtEqtRZ
RCJdZVYtroEoUg/po8oUMMgRlcsaZgCq4qRATPLAEx1iXFGHVqA2PHjwAtu0ii5pXAxMK2lM+b5Z
tlOB1fNiaKI6hB8zuCfxuugnbRtjFBWH3I6AQHducHe4EB/r4miB87bGHJgDPMg1otl41u3+mOOn
GUKeMtdReypLke+kuHgY+qeW8SWdJuQBlAVHNNb769F92IE/XqPV6rV8PrzvESqmvAQ4OLOOh+gy
JyN7WL6B55AckLfH8VYE5r3oQ/NT8UJfN83g+seIbdwL/eLD6DzuhGxVMAMpqltgTIc5jmXme5Nu
Os59IommeRmXx5/rAXp/w7vIBj46XfFtzcC2DUC/VTZqM9usPOO06bj2G5HyTJskSceviOxSPbKu
dA94pcTd+Id0scdknBiOtNUvDUsLsEA1IKzNELtEzgIW3nLbEsKCywNvbTggnZ4mwDG/HEysJrHT
l6SDEgasy5ZjSEyDHQvgiW+XIXFfJesJAPt3HaP3gwiQOlGen/qRnp1xJk3wo80s4YSbckvRCsBr
Zk6LavLkBZJEqb8BGqhrS7RaJNUeO8hGu+ZdISZydLjQbaqp6lhJASdd6FUNVFWm7CQGAHa6MH7F
SgQX0B72I8DJM8Ayd5Rm8AvG/6cmO5fykYZc6gZyuN9wAbXIgynfF4n9EYgG4shLPpP0nYkFJjsx
0GeBYyCwrSUJ9YZz1pDqXQpKSQV6sStUFVU2bfz2l6QSdfTvKQJ17bE9eNvJosPvHyTJ0tMhMz2c
m5Zm71MzF6jdJ/yR8zUwivZGyFrH6MG8nJNTIr/1eP9JriWId1utczKmBjI6bi6NWaeKN0wW5RTw
uxKZ/l8S1+mACbuX+4O7PazlLFQ/b9xda1hiYt7wB6sUZthtZRoWsGbB9rpTVky1GLPMHd+Mv2B5
9eN8iYSldMQn9hvJzYlTaH862uZYQzy2HNIIDdT5K9OOhjCAXduoke/PDNCL0AChSwI5GOQUu0BW
b3nrLfrULfIPmurFUhsVcdbf8BbN9ChFKnpK1j46gmYxwORMd2XHGwZvOE16+89D0uApzG0JmESh
gqiuxH2HYyvAnKIxAl00ZJ6qjENl8dzE+KhfkJDJI1XMPPov/kp1Uj3ijjCBo4lgwAZHs+bTXR4B
4NzNZTHoRP+N/+8rR3uy9W882xDsalfUUTCCIO7NxixwfcnP/DKCpitFb2KPVoUMgkevHnR7WCI1
gArG0kLz5dOPOvO0LwZqh0HrpJ+SAzNNmEk8dJbqoQ0NG6tmS5uXAS8OMlYPNTBTTrGWu+NXcNOo
ImmUNQ/+5tSv9/d3YParGphXjx8YSvAt4dQqw7IzO22fy9kDOreMMyjMlvM7tludDGVVcgM8CF2P
TuDEyYHwRbuFsVKrz1MsRujubcloRi51IB66nvc5fu66KI34tEj7DzCICxqDj2kJmlRMeqAy4+M0
23qVtWzVJS8Ob6kep0cc+iBKk+GrUgN9kk2Li5NixJxRNhBt26zaWUUsSaEbwHpZKaF+xAbO8sCq
SfjRx8f4JuBv1eD8sFRJC4yiA8mdSkR/s7WnDdDs7fflYxCm5QT0mOQHQ5ZV6+XXndwjzbZ4FIdA
dxdgjRojp3/oYRrBeZ0khwm9w2A5IZ7RO+9lTpC8Frb9E/eQdApBeQU/Abrpg9g2Ad9aJvl4BCuF
ETtm29sX34V1s0Wlw3f2hnITSvUjRWNa7b8VIYIH3myJwzfilbFkArspu8kTSHb9fMCFjPLZzl2j
I107h7FId9r4eInLERmGYQyFF8eWcogPR7E16vcMP2fJi69V/vFi9kOKAcTqxOKH679Ef4AxQugC
4cd3NXBuAiO6U0NmupkqYcCq0c5NTWSR0PJ/jeOerpD8VC/1YAPSfvv1OusbZ8qe1rXJcSsuDPBa
6uxI4NR8QD9fPVVeqGTyiEIh78OTqWV9efBcWK1HxjtFslOhwNFkJMsxLoi86RPU6sEeJDpR1Eqz
xkOJA2rIQ1yiwrRdPYtWF3X/zv9PE3fKBl2Xi2W94uWHpdBFcNneNPfgC2iF6JLWIXl+SIgCGyS9
NGkBW3+257EnFioi9JrN5e0DUIUMcI29An1OUWGyEKbg1JZSdD1vBTL7l6xMS+pnQiyX4NwjitBP
hARpCY4UuA3a9jdzG3ZCzHYc9TgclvHcdfEaEI4L+46o59hFv04uUhK712eZiGqRN/7wzkRKbeHq
eGUXyapY/R/sqMOsiNef5OMVb4CrR4fcl2+ZORaFpX82InYbrlSmC8fytMk4jVKPag6CIS5KXRvv
6EMfGHD9YBlPneC8Xp3VDz/T9QnYEl/f3mlu09p1rxKNqgVxWKe19OWCv/zOHTHKHDJqm94GAbBm
Srw+R49w7Bh27lcJaQ/we6DofLMltcSREGHjEI8/rqHRpF/gABmF3B+0Lbxz1RyNOzdAoUKRFYPF
Fwzj+o6AeBmk9VWpTszqKVDo/FAtBKenCb1j8fNfnW2jjh1h7khicWo9ZHVnul99a08gLw4u940+
N6UAlhKXGUFdP6pQGQYIsTRvmABuDMU2rE7OZR1oAy0fM7UOlSD+oH9d7e3uzdwcYssohuifrSSG
6KW6TET3BkZXpN3T5ATYRv2R4mnbzVPu5PGRVHLdF5XfRJi1evNIE9ZVmv31riiawWLJGOLEQqNE
EkBadm7FQajzJB8lLyMj90N5WkqtCEwYPJpHSHwDBADqfLl3gIraAbROQhMpJHUwJ3RcSAzJx/sk
tDbCYI17PyII/JcacBy90fxhzVCV4ypO1VbWY6bHyA44c/DuTGM91aHYAjujgmXJzMSvb5fFvpZQ
eo22LxJs4nG2LflJyQcjCBT5lHXZmm+grSuysMNzTWqJmgZaiimpHgnClmwPn/Ec5Um5bRy7NWbV
XTFhqADDukTn2r2SX0TiueXe8FyJ/MJEkg+xBsOOxTyB7ySvV9EjtKsNsCq79146po1lGEJvYXNL
vQ52nupzmWO+8y+EEqY2WMMOQ/Bj7ot524zJHKvJ12QpcOBSVbhSB38YJuQKzw1kXMxC0QhhUisP
IFfj9ZCY6VArevkoxzWz5E8HXX0yIuN7cVGSao201nD4xOZQEpfoy23nf5P8UX4hEmlCxyPTinef
vB75SU/EiWWdxMGtQ61rroc+83/YPZI6LWIxAi2YPGU8TBPQvCSrZrcz9uyRz5m0yE0/m+txWhSM
yrVU+pnBxzX4T2lpjGQ/ZuZ96QgdMCaeFRmjKQ/J/9SitoOo01Jpg9cXGle0P+Ig0qaRURjRX9Xc
uzoKXOQlNt8SmeWEKQcN3YUbpSEF7pes6zVXeD4bACVu5KBXp1YiXBSAqn8lJZ5p2ci47ESe++mW
1H0byfzeE4cQtO8TrDIq9d6oOzKEJo/rSRwq1VQmNgQZPKrBAa+R/WTFMXRnK8d/++ivQJetbsZh
HGiY+BkI86MPfSd2xf/B5I9Rzk82ToT4OMoY51i5SknU3Ht7lFvNxrBZakzxcwV8R0wDpps0MwTD
zch+y4MIMEeKrTP2oqNs+GKTxgPPq75QbkVMErIWMX2vEx9SGDJsIOUnIN1fj/NuSSp4Z65dtZJV
2JTA/sdZGqP5Wwzia2ao90fSqYZpxIKul8YZnwi7Iv/8dZ/bmUN2NDPzN7P3mVPS2juJ667fyB7V
Cqx0IJvaGrzoMmUsAmj7SMvji98b0jlI+NmVRpGqdk/H53NhnFhB4FjXFeK2XwlYKp9BYQnu1chh
BmZfUmg4bBB3DCoosjcw0Ery/kXgNx3wPpeeZywUXwPDasA9J2Ol9f34AZslZcrMg/DtWCIN/nsB
6BccjLBup6jEjjCT41j38E+wn7DVUDpx6BieJnKJ/OhUFO77pv4VRk+0RNCKxQDeyGfpjFVYnzrB
QlCGIchECaHkc8WaNLJV2M3X7Q30L1626rQCC96e7VNoi81adSYyd01tCw7k8ju/8YMrbtcxlSfA
sbcUx3GsiwIuaw0eO5VV+/9Ha2Hqtb982SWwhMdyzORXph0A0YvHxnn457Yp35SkIy4x8fpoJKXu
X4gRiaS9qRKa1C1zixiBOLMq1+yK0HjOmORwwYQLc+SKJ7gHhwqlTLqnRSYodf4N9dc8MEAF3/mz
3yySOer0kzq0LjCwdSIcA9XaFy/QZ3ieOmc6/SDB4Ib3GDx2N9vyUyGrgBjM4lly7WeYy5HlOFq+
NGWm7Jg5+b8fimSORAnZa+1R9wQZ/tqi4eMAJca5/gWGltrTmggAgPrdzzlpYZHejdDqjLT5Q71M
BJ+6HToYBTXCOFgYYXRsgxkv1z6ywZFS55nsjl56Jn+kapB50iBQO+R7+seulc2VlCdxw5q84N4m
9fkPdaOhmoZb+9tmUqhXQJrS21TizOuEv+QkoKq4dE2NHav2Npu41ZXF0tlzJhnV2wphzDh6CXXb
YpMCIiIYUF/mllw4Yf2CTW2prp1PAmk4WfQHo7g5xaMC5183kUPTeHD3OiX+N+L+03bCN4CoepVz
GdQxctQqzey99lIfa5pfJxehbbQY/m8o+xQlWDdaAq4VRGh/UtpL4sPNA9dJ/yeQQcOGMFnrz4X9
XgE2JMPLg5GJh3RrWDdgotzGjbauMv9gEEmKRuItKiJQItWSQgwPDlwY0jZtaOs45SoUVFYWb2GM
UIXs9GGul34E4XaxSaZSzDU59aOKizWbayOrZADdKwqCjMIRb4QfV5iVWskNFD5XpFowLAgWi7cW
PrssjKcxxpPz0+oDAypmQ6x2idw7RoWhVaf8fc42KcngPieY7R66cJYmpbFTUvwTcXbRGiOSG8l+
ZlTUq2lRNLJR9GgMXwSM/L8PcT1IGB1qhEpr3xDnvbsJqPcA86KBRuFom4WUA4TQU9TW6so0OpTp
epEr68N4TdgXtOYiCDQqHihdYXCQ+XDYbiHoGmnsR/sdzT9STH1FwFVhg3r6ox1mf4a5SItFbw7A
n8BsJ9174yPydbbneR3Y7M4IzrWaNuBVn0cMyFQfYCgRyUQLLnXgFS/tc/ltu0wVov/vMxlTqKyD
PQdcm2hcKgYlI/oygLUtk8qqkBTPncUkm1L3k5t/Ak702oe5k6CjJ1OD2lUufO88jbsSmwb26zNf
uIbnnFQC8bOVF5A5dBbD7fjda6SH3dV3nAvnhnMCoqYTY08khW5oL+aWLFBv4+ya2H6Gu/mMQ08V
Ob9cch+AjTSE8wtyy8tiXRck9utVaoJOG7dzMR/ZT6P3gb9/opVYe1Rtnt0YHH0O+t0u6pZi6Xo5
hZ9eQ/bCaR8wXi2EMFcziprlZiPHcH9iD958SsSG54PRcWM0hrVN+2zh9mdfDmnjQvDWGbbSlZ3h
J+KHd1d7ERQgcQ45uNiWWAPk1UOUSEBFfN9EJOg+O3ZdcsMgU2/q3tweN6XUTYpp8XGv+1Ty15Us
RbR91hAjpW4yAom0V38pJkaoDcc3LTWZM2/nhHUcBba8dDmCPgoGEI7dQzoKnHcXJpPjcQe3TT4t
lKO1Fba759bDQWKsXvXkzbN7DWNLUgBD2fxDs6sy7SRN/8Ep57ByeElIJaO1NpejCa2swZcmZwj2
QU9jLVNs9Qo2kiWYex5yORUEOZ3DLvjuLz9TD9S0SIHvAwJ5kYHqh0msjOIs+4+NwbYy1CWIMf6v
pYxADFex+rloQ5AGW5CgJO2yWussGx3XdzAmXNZT5iFirOVZ4v3BPBy1E+nDBUEC3KJQjk/IUgvf
ys8UW73B6TusHHIrBakq4YatKmOAady1jjgpIupK8QIdF/+3TTM1iFvMjsHWHBExrnPqmNOeB2o1
fmz+qJrYCQzN2U18P5rSmUW2vsJ7wRcpEKGipqQn4dIQJJqGIW6zBngBPCkd+HhVSBO6ewrF/h4v
ad0iCHZfDrEQBBrFtd46Sw1mSD3dWqo8v4JNMxNVH5g3eLzeqStjN7l0X+lP2Wo7lMLuGND8yWLq
GW60WYUIG0ZIJ29AuxSIHE5Kum96HhElnwSax1iph09GjbhtocvU87OEpmZSZ+a4ziEY5M+PvZ1i
dmXzjCKcooFRGUMzvCy5okIAmaF/OhTwlvl7K4GWxfg3YbR20rVejx5ez7+LotSebyVxtbpAdtAh
6TbMq7KTXzAe8ZdAzNBGBBZ2NXMECF2KGmZuND2ianBpS+GQrTOUMCxrLiTrtAw+OnY8aO5q+H3X
VNc5oM/jgq88kVcNM3BPwvvaYJ86fASZkwFot1LcyW/Bv5WtyTFtbgiI0A3CaxmyxWkNkJ6Xmnfy
ArsjUHbtmE9eZWdBCBMsJ1ftEtgRK3Jq6WFXv36ENQMpENlYzX5/zhZTeTA9O8b6JUv2a9WjEvGw
X/d6aZpOrRSgIlx1JD6aLtNjTy4qM4QvJ9Xus+4ld201PBc65obw9XGMJZcJUybLAwBY6t5r9mRp
cuF5RZvsJaHO+TOYUDg6jV7zMjeJEojEFRqnRXWkaWbkRuyMuDXMD43nmiz35sNfuxYithmGuidN
s1gOIerEu8otEnozeHu76/pPhYViLmO0OEkf9b743EYiV5ZTXmUtJIdWbutagQpRFt95fyUXEZGD
f23jd2uz3DdA9zyS/6aFE+OhKCJ9bY0zDHCXyq5vD+DQkfZgnVx/3yfmSAlXponh8I24PuhjRVjZ
/8PF2WwYQmaamviJu79paOus0Tur0b4hWIg+Dik46uFp1sDxGD6yp5RyUmM3yhEaTTMRKTLVnlP4
4zQ/cBbTuKQ4dU1TYpYhWufSkwNQA/pXEvTAcjLMaYpYhANHeZ/h2E1NdHCzA/VhxaQEuTDLI7o2
etDCJpn884T0xU2jJXP06c5lNbaeWTwJm2K3WscQZAxLPe+DgiTnmbtdmZvxQRLSi3757K9VFfeT
AtM/5X43D/TKf2ptuQVU9iKhHkzUUtW0OGHFX6N5D4Uv0u6V/MKCNVYniKZ7nrEupMaEaIh2REY2
BGHKMDQ4lLxPRsuQM9vRo39nZGJ+F6Q/GAvg7LCebSzhhr5P+GnFxjV4IOcYO2ToEiYNh6UowHuJ
MnRTMFomivakgvOiF73g5Tny67ZZKX4oNYA/vMiowatOwRvotC2wv741DcPASO0KnA+5UAfWnogr
+zmoazr0uji0Irt61rUd6wJntvGm/HUJkPsn3yTX8JEREE4QR5jl9p57cB7Xlge7RYZL4Np2COu1
Fccg0LWMhadXayeqv2sC99QsygtD+YeHO+MM+TefkCpgvqkbr4RVLQ3TNDpgzYqfh2Qzhs8R9dj/
Pm4MrSHj7onREuQk+v9vRLM5ioaD2R24SEYhBscEXdmtOiQpr6eXFKnowJWrvHnIGuGo6i5sdO8n
ICEJQS9BVLz1qfa1Xgco6sdanb0yJLZssWDfJtk7LsaXy+zIXd9wSWU/0Oek8YWO7AXi1QRh4R4W
Nk1PJzzPglx94loExZ1fjyh/1auDSS68tU0lp5S/+/2//GK/fe0irgN+oYL16BnUaPE8OftdEtD+
kn7Er4KQY+M7/m59HYL5P1nHOI5ycrSo/WISkKYYf1sUHx6JWokq30s40SaTOYdQrtn5DONkPErV
bJcL1ldwvKR0IqJmi6S6o9OdX2Y8lYEW6UJidQz0Hd2mAdrFPXDkv4DbwMqQ9IBi+wM4XAcm60Od
QK3aB3JZL9kUklAJvm+0Xw88vz/1sRUjZeVwpLXricN1bV8OrbM9mA422L7fuoN2y9WHb1nwv6KP
l5M4LqcXFo7s4fHyEjwbMyrenC9pTG9B62lRyOy2PFJpwdPAVm60wT/ud54t8IdNkknVOp03tgDb
a91bANgmhDTmvkHrkmwEO6twRm58rmDftpCKocZBS0/Vq3wgMotCvY8HDAVdon56KQXZAZt1kbHe
emjhNs3ucV3hMyRmvjedmNGkQRbcMheIADmlW5XNsDHe6ei/XkiZ1akVJmv3oUztyciNraOxx7Op
G93CVWd4CZt63qg1MQ9jW18a2IMXQFzmI2piaCty8Kpktk5Ahoi9wDTRvd4cZeRtNlbAqIEnwafq
XELhUgXPFbcruep2f/wCCh95ohhJhY3fqO5PcCUjID1+rJB1MWURIaX9tBEvDgf5X4ega6c3uXWB
eZDBN6qfZHqGZWnypfjfuyz7cuaACfHx1CRAQoCK67T35MseOrmG0UPqI24voyUvcrSa2LWnslkh
SFYVzVsVg6y/jpn+GqUyCjeLghUMYZGQfcaU+L8Soc6+gYqwYyY3Nxw1w058tOg/R+cTLycIxeHI
ZFU4SuvZOEoiR/s05kpzFjOtd99DzqngVGiG1Mcw6JA07mfG5acYlGvSy+td+sBC2cxVtNHQmV0N
mcyuvLMGeAhbBlIWHSzAaZOG3ShwAWu2uxvxNX5ex/hrsmEhLqScsNje+F7RcIjtSGoCl2vm8/mC
Q0FGY+bIvfbkHbnFq+jnxoaF9hi+auZyds/HsusNOiLlAVbfrOt3DbZ/OKz9EvUAsyTpV6Cfo5ym
rqYSsIsCYKCiA90UE7DlrNVb969FzhvpzVBwKC2HcAsjWy2sMrqP46CLqoeDhsAPFgVmF+cKM0Xb
1aHdXfdrwhA7Zot2HmqF+mdL4CMVIY+taPq8f803KxWBzSFQqgw8xDnnmuibehw8WTwr1oxidJpY
YltrPjylEm4cz38xDnHIA79x/I1rGKnMaFIxG05MciTGamb5Ap/529ZNe8n7SZRomy40nw7RiYxb
0rgwbQCOYEVXx8KNd/aJv909xdlIxf2P+D6S2NEcOyrJghqAa3GJkc65E8AqQApxwpfUVmo3ccZ1
B1zYRG2c/S5E4RJD5A/vgCD2IP6zSHLMceYDKefLt04NaFBPi2BcyczXcEqi4oaE7tP07m/J3tGo
Vu6pPWKkpCb/sFYGeoICjGLUI34M8FRpgqYRnhL7nCizIC4sC04/2J1BO0DK/mRQMMtbdZdErlI9
BzksSgInpyKC6me+dTwFxjYMAEmAa6zQ6Di22k/ZiDBLOoGLF4WVc22a/rAfKhx+2f1VxR2xf1wv
pThaXTk3croE7q+FaghI3WF9B9/5zjtewVW/ybdCAqH2lmgsIbyuOCjXeaiSv+KIQfsItm5aNRlu
OYgf9Ed0xFHJPH+EoggS4wxL82c0AwPFU6nH4WRugH3k75/A1sX+8l+aNKPr2bncXkryN6RQwZUj
DP5yEDlkoA2VhNU+QtxuIH6CJ9xEcUJCoJQf+U0UTxihoPBU2HUNt5DOSRUbrcip66pM8jfAxrUu
/g48EEcu/SNtkgHfe3DJJ7H6rAEzhLFYhVn1Y1AmK/zgDX8LyfcejuVbFO8caNzUCMWK6wGesWDu
4GbjYH7ldfGIMXNMnTzVH14T+ZntxFFwoTORg23i/1dN+zwgRc5nEAstp3of210Un8boS3CEJSkG
jBZpSkk/F6M93DuLahxTboI/MwDXA+E3QabsuMU5y04jEv/aV6gSC/x1E5wAE1gEkWsMs6TvH3EO
xBHDPI+wFk+0KXGbU3ldQdaSS0cPU7+YBIvD/VXttp5W5QhSduOp3giKB6zyZzsSk0qbOb/GYfTG
JlwdsCleQocddGZE81g6cJfDJY1pv3BCMX56wu5dypvhXX5nmuHxIsnPWyoSuO/Y3wfar1YjhHUC
fb5nNK6C+Fy0vWudI76QrzEq8tbvokWMXU0EdZjd3Y60xZ4af9UjEgGaODiC3i+ztvcqn3g+wkuY
dgpU5/zRzzBuGi/HMkVOhHgwVJghv7gICrCferH+P8DA/FePxd45bPDa/JGu8gNYn+gRk+JU/fGg
iP1ughV8vja+ZrNgLLtAscFbZwrzkG0BpmPvDTrkuDQm2I8N9Vq26zH7TwQiog00v5e1ICXjCAkK
zO9lejlWUuKBANGXHcRVPLJYcnWqXwCGBi7p84YMKGAcgGdQmlYPtDNxao9CKVQ6xIWCsppn7NB9
WKFIPjEI0Al007JnOEKcCp/AYfq6ZY8aUQEtJRyiBqMgrlVgGLgp4Nfb3j4F1+9mtKFCr1Jk3E1g
NroXKlQostb1T5lZSMfp6LMPh7c7cV9sEBshLFaP0AUYzGPE1/9Oengt/4fczhAjn3V0cg/bSadt
8J8YaRZNdqtFB/80CpB0AMNSqjcO5X64b0+59HrHqEPI5lYRJr4HDC/oan4lkD5c/9ybplWNgA3o
MhW3p+lW14pOVi2ESB+55Np84guuD2b0NnCcVPUfP21j3bQfeZJTVETYuS0/xe3pydTTote9jww4
LROx8LwMSpYMfjWcHQZaPXCiykwaE/Vj4A3UXh/tTY93fp9S1MeZxyN9XbS6zcrd9SDWVznLc/xj
GuXvGhO49QFJ57HBOab8svRZbw903bw++o6SeBPVueqVdyO/W1Rc3QEF3p/eidixP9H+JTaA60js
aLPCgmnZbs0P+tTR/1mnK7US6jYlVjge9O/rGQkZ2JFXs0vSnjFehF324mkYv2WAtIHmZsouYPVd
oZBnEYU79ekm1UVsPCxwMoD0I4LzTV5bXsbrqTN0C5djUUxq4L4qKy3oBVzhvFwJQkWEFTnVLTy0
b3yhf0oLNTFw+dV37oWcHQuPo+UNsjS50XIK0V8zKP0x1u9Cqs/VfrhJivN+L+8mdfhrAorwRfuD
ft9DKMF7TXOPe0evrZZOD+Gxuz1/gaFeHT7QPo1obIht3zhmYvk5oED3XE51c69gTs4ZTuozvsLh
8oy0OSeI0pvgWGuEbEOMlwAIBNweOMhTRhR3BJlfh5obR/yS2BCGAm3Mhlf3P7taOxgLhuwb+rv4
rUI3ipIkxSUS7Pq6Z5yCDA2coRFURXJ4lhSVsmpxqmtaotoBIZV3cF6imRsY70W8CJr8cSlSgNui
3AF/2DQ/vGbZ5gyyuFZiIqOfHcKElP8NLwF3MN6rRRKwkP2VvjaaRjCToa5ldtrFF6rSZTGDTYqD
uVNsiQuo9qQ4X0pmGX71nMtJww/gu6PwRAzQ7MYSJN1CZ0zvUSRXc9fSfh/VSZSFSLqMjfnmNbS4
wSlVxzGd91RxnIjWYVovVLueP3HsaDy3+DjEzNZXYileKHJZDfwHPLTpzLvmoIKCXDjYmx9Fq887
8gZodlsBF1ToX45oSDfVilm9yXs3wmIBSXU+azddjb/k7n7hcvYE8unHCMxdB04l8ENY9Y3kigTF
3PY7tfAAODU4s8oN3uxwMVcd4D4WD2P0xuxkcOdxUqoLu924g1XIuHgICgNfl2JDxXiETi0m4CuK
2YrzbN1o7BX9puNp2iv4bdB5i6K1Dx1JfrRbNrQZMliG3Gb026hPP6bgQx+ZquajCOPt+XBlCTS+
w/wP7fJiRjLuxGuNy24HjaedO0XacSD0LXurkvd9F3QkNLEli9sidJe/60P/10HE1UVPg+lyW7tp
FfPv9S3ihdM6+HtkM+iOwBBlfIejzT70fG/k5MxUadYACesU6ZakdldqKsXnit7UBI3f9ySSMvzB
DUG161u1/tPCCO88k26kGaV2bcwEy//ZsxZvdl4l0MsL6LUHUh6+1tT6LRb0Is3dfN5VltRxUfca
5XfLuPhZ/YLzGy5RZU5358DMDUZrTvKPvZT8rZflzWCTn0SfOLV0UgIPEFytttuvgHYmp+sjzihp
apVDZ+TqGODsVBqXT8626UdX2eyhAhbz0YRJPcXJkiIMNS2e8dSiuboZznj7W6IyZdzPR3G6Hajs
fGEheqfXYj3KBzH5qtZ1d9CW/RkKDDZRK8nJ6drvZFH6Sl+6AKADLd12e+jqoTSQDUl7/v2mQKFF
VJRQQ88rXkPCp9zPTLEgYHI96vjXDCfjnuPDIncQjhJm7mv7rrZeF2cDnpGODFu73pXXc2epckNy
cXrLW9gqoh4XQkzSwy1kV8K1PjiGzM3NOJsNul8zqF6S/zNSm8NFmgEpFhtsAqBjw742gRr4bPdw
tZM7vWFaMy86YWJEsU3pdgQ+dLan9+PBe5/89M+LYC+zW5UO3BtZnSnrsaunC1rFUe0tKmo7dnHd
liQspLLNrFAqV25mwrr27YAvaMby80pStPFyWPEhh3KdUlDbBlVeQccTaRcVux+AB73IMA1AFl0b
ydKuyWD38KznTRW6nyEb2RhBJKb0eE6rVXSO571pb3D9G/qgqkIOYixV5M6N8YOwoMCc9HfkL1r7
uoVG2lTvcHkRuBDlC9NxayWbW3wNOgpu1YbNk+BI34vz5Z4Gg1C+jATvhsiUelg1E6mH/7FV4Fft
KQ+wqNWDW6WLX8UwTtoK6sUP+GbKJhm9ujj0u7lCfSh5annI1UclwoZdTSM2nFEFwOaJpnmAFv4g
jxVS8rpHnhADtLLY92yn8VHHyDOGrrebT4+lGYJ9n6vj9d9MeGxIYb7CMHhd0GEHw0Iu1O9nkcXT
9zA7f/dVRQDmfE64KVNY8POlczzm4e2pTh+ghJT2GerTuxMm/FyFgFRr7z2tItzIRiExqFz25bPe
pKbc4ufQ1xd5av1oE9x002j0opcSPhgbXdvuNLGqmvBWjll4WmBO/vR/T+Bz5mtl+eTN52y+TGIp
ATxgiDf59a2QliJCRU5i0fbhDEusGTaCwLsjnHEmzXDfIiH0ABQE39FmlOAnyvjOSoUCr6llZUsZ
ZNkasNLgpref/2NjycKfUfOlPIbc+bZ2TNhU4X8GWT+xqvRPxlOi8gsyaShBpkiPcIVbYdChOB6D
vyW4AQz3rf+k4ENFhqWjPyDFURMcg4fbuo0l1JaDuxdSjiQi1BPDuJJEgZAUo6Z5NUHELcXJ/f16
6M44/Ik2h+r142WTpsveoiFPm6bujvawIoTYWKSK0WqncvNPxuCCnQ5pG0ucsTcBUP57ou3H0WAa
8pSate8o/+p2zO2CQqV91fLQny1XqZFh/+Tyt+VKUf+Wl9JWIjEwpFMxMnQJAF85Sm5509WrGPS9
iBn+nDZYiy8HRNfc7AdsXDoBKUz/OYoPgF71FZ7QZSGWhcvFYitG5PfDwr8M/sQ+WLpM5ApjfmeE
YnDJM0ha5K1Q2P9kLMIGUFqYTSRXGnDL9GSHhuRimBRtbElnK3np9/jlL2IAtgbVws33JEZaS7ND
h2/S/QSAtyPLSsOhOIKhEMZTYBeBB5TuiJDhNi2qrFwUTS2+6NUbyWo07jEQFzHedtdsFOjZ8K0S
S8YHB+6zk2ba38cvWdysljLLWckn8y3hJg339banmrPGP8q5nIXpfVjGg/AN3JBFpJf+1ER2u7Fr
CZnaDnkL0IccPyb7y2QMJ0ooVpnk2sdYpp3UFTJ3epgOCS7SBgWdc3NTHBKgY7h2YFnLuJRKqofx
aQJBrJmiyRil/mhOIU1C9PGVGHf65MhrtZMqFIDxCWe3+XZcSTxQ+Zoq4wdRr3x75b6g4M/X91pO
kJzroNLG0Jpn8B+z54Ss6VaL7npq+CUjZN2fh7qpw7hmm8epUT9FmuvHTDjtiUDv5z+11IJ6bPpg
maLqpRXe1n2O6aoAjEagDcliJW+ikwFcCi5UU2bfYVLijgK1SywfBalcNFZImRrnfvJHcLQ/VkPF
njea4x0Orn5+D8gi3HjXadIGNrslHnOqQ1GmHvcl15+DKC+WgD0UplxDktYpCR6OG+65/P28P57x
GKpcbBA9vvCOIERmq1s6nv2zXWEzlXLiydnRi1c5J5u+0aRgvXVxdwS1m9NeJB12pHbyjdZ8R0N6
9Jc5WMxjkHmgxL7Z0Q07C0HNA8YBi2AhIYaDgTIoAHUYacT6Rn4pX0g3mhTDQCDTItRoFf8BJzVW
fO19LEDEwI6THh98Dq9Rizkw8jdDfmwV2lVlx9CIV782HX7lgmYijgirIBL6LDvz08mm4qqYMZyP
0CqTEIVc3rsMcnD29FZi0FGf1D3YB/TvI1TLW68NgnRGXOuQZjrwFCJ4s3cXECPaPFAJbSfW7NM7
0+nJXOhECufMOvpm0POCvUBqrIARnZ5I/dWm4DjV+1uzoSIP7GEkO305NERma5+7OJNmTdcgZBEK
X0EceBH+hMPqnPkOCKO1D64D9PzZsG5zQT68c6dH388MqDH5izKxy4o4Vmx1j1gw9FAouCGZG/ir
cjSzp0EUTSDWPSYDZNqxUvqx+1IrCjdQVSfiCye7H/9mCq0qY6eo0U2oFArk/x+fywvAkZS+fAsP
mNyIR3SSfjfyCXNJ5LAYL3Ac6vQOa7LCKBcKh+zBw88HaFHOgexQlf5tR7sH0X8DwhxlT32+n371
w7Q82q30puKC/kRlZK7eQwjYT9CxiXRC2euoQpWbk9tA/4RLqaQN0I/WlXu18JsQeQ8loSC305Se
DDsp1J6iNG9GbUznLbsjy4PeiP/XoU/Dl8w28+hTu4UKag0rZ00cQKYXDy5TiWqJqj/5n13JK5hy
ySy9JBH4j5IFzMM2I0aQXBaFOJgRe5wrynoTWiTOb7+kVlFA9k7uudRQreoZjQyvJ3kgXMlbS8jp
qO4WvG6ypatE0El/R6PfI76JSdFdmV33xc4ZJG0lO1whtsghA4MNmNRKKUnpq6YMzeR3xvK8oipT
D5yitzTmwEbVtAbWeaItutzQh63NaVD1VRAnGmHKeUfMDgJlfNuQdbAdpX2YPPE8q/0su/fSAglu
gjQvBUkB8gV7K2KrnTnRXGmsnex8JZCddP+t6qlUhmTjSp1Ihkf2x3Zpk+rK2uPPGDqhciJupRdq
drTAfvPwv9ZiSfGCX6yBM4X3gkHrrl50iBXGkcOvsdas+D+hgwJAarNvTcBL/j1CMSjaj6L+e+N7
tokUtOCWQoOmyV8PPhURigX40lQJZzQ4DSfCT6WwaUCpwAc9B6kGOe4lIIj/lUg7m0ydaZo7WDld
5B7Yfo8OLmgPQAEO5KZw/yXSZzQQpcUluhdBKtwGvmi+IF73KmXjBfvcn7RsPsUENjOrkzq4wmUB
QWUqgqq7pvoIBzfQ1178tTuZTXqKSXx/NDtfaqyQ0x/YAmjz9Os/UgGkqhx1dk6/WsGa3MeJ/4V1
ty6ZYjS/ODX5RfyVfAv/oo6XGkDtrAG54RNWJaHXKGl9Fqg9gs03bx0lZHB05mhFkJzzv+JUjfQ3
XZYWyyxttD71r4vhXrWULXs6rMOxiPlrOkR8PS4KrmoZb0XA1hhT88MIv8ay4aQJU3xxI8mXfoIl
F4WwDFgc0md4JqY2Z5JlxTeX82nxhp4PXcFYWfJF36Nes5PonpT60j2kq8C64jOTNLitck7FvRbW
M1WkxU03/+NTfw2VNZ0NwdqGtiMAu6XTbcIW7ItcYzy22BOQuxfD2pemGBNlYQ6oYcXZ4jAAmpq2
jJqo1XxGrHc3cMlg8eQwUa0S8JppEJ6e6YKIFgptA5U1ffPQzgQjNJlCSIKk/6AdkeLLCd0hn/qI
3qx2KsDSCD7V6V04UhmUXkuW1j3J9ygZmYIZstDx9kQb1wdxaLtw845Pd2e96lBEuKZ6WsnEQjP1
8yx1OljVgnjbWJqYsm/UZKDV/yluddyan8fwMewirFrfeo26HFioxH3xKLR9Bq0Bho0k+DfLf0bc
OpAmJW/wio9okY/art5XNlpMHwz/tM1pzlrwYgbsm979wpjV6+GTf3oBs4RcJ0NrwSvieXKv7RqX
FxwFItZwFCkz20r1j90+KAs3v/d5iibCdrW29RNW50YX0qig3/O0JQLNrQXUmfSrSAJAv2oq5O+j
+xTfvJRzUsTFozkDCsAFexQJdbne+Zbh2EcTbkqoYs3u+0YgZZfnnCxZe5TTG6bXhnuT0Yt0wjFo
gssXZCqCSqY5WwLThQBIt9KGG/AADn3oWRMUFU9UQ+K8nreI5YITFCNRXZPoHPoRMLC1vDIARWkV
7MjnKZk38D83Xg0w7XcZbSoujgGSJUDt2FO+M1PYdYXR5J8+Y8Ggs1WieRpjjA4QEgPintAHpVBC
NnadCNuSlAOw1GEzDN3e7XrSYoQmme424dYbseW2pN3YWR1sTDFf/RQYjNba48PN2cq36WUNPlqh
nmj2ZsjVld8HgCnWnlr5EQVC6T9dyBpNSnJJKNM3uFUf0EXSSAWjgYJLoNrmmrDNPuRqR+5MpQXW
04Z8kwRp0pM4kDFPARUPuAIjMPJYUPCeC/KoBoP+aCcK70SWzYDWpsIqVZ0GdVHJii/m1sEJhKvW
JOfWw4lc7spUR9UJ+SgyjHozhHkstD5gZuztI6gx/ZqFomrwOzRZLvAiN72aILAltKGKrnASeYAO
tEHQotz+c5b8e/OExXNTwLz2Y9YwNOk9M67eMyDq0vphN56y/ZEkvgoqvQSJHkn5U/l3OriwPiAR
KcqiuUcMDz5sgiXKGoCivNiCMKWCpbbGvWNUu1H9RNs9r4SXmIhrRDD2tRv3dDe3DHUGfKE/r+tA
6ur7TVnJZhP8UL/UzO9qCvXJcqn8+wNQZVKU3TGhSd0F4jtzUw3PME6olmWdNRLBUMJaiq9Ts5q6
8pZQUEEcKOFZyEV+gENMX+0KMzrrc3TqbuaTYvWkjrapG5tcqGG7heqh4fzjW0JJrFHama6MvZ3n
hsaEHndnfTAKd/dvU8i1IJyYFjaH/mtgtRhEGudY5iqr1E3tLyHNx9LYqqHOlyFv8DraAI2AY74A
0tlWpUtYWif6gPfT4wpQIRkUUSlBABsaXKs1wS79laTrITWlFU2ojoOCD+PkGfTCldYYgG5Q+NlF
/3GbI7MkCtr2h/xg8dkd5YbHfq99koJ5Tp2kDVQcGM1YMFNv5NikwrxnPkB3XkiaHwiZZn0S+FY9
UXM5A0nwSFW+0vvYHndIL2AwTK88m7RUEYV+9NwCR8uo2Bt6kpblhfhWoOzJdoA1627E5fJhR5Kl
88NrdEMLfQGkOPo3/XY867InkHnmK1xO+Hqusf/vOx8s0FyKpastVevtuQzWts2prJbjWrE2O/Ka
lqXWPNTZDfA1OfYieEByFXfyPmfilTZapQrTweqpgouDArLjRp6tqZtWGV5y04TXKtU6PGhmGuqr
M5gTz3yypSxGolvJP3snt0cGflgwEt20cBX/8dmBY0n3pic01pAJ1o6CDxyQEgviewPE+bkB+3Nf
SySwRjopIOVAcBct5vTnzukX9H3kuBA3m0VaOq3rPOQKnS4M8GG6rNyw25cRHPfC3fOCJFFpCMCx
+wvz0B1Zjv8HxnFv4jhmHqM9kTcechaI6cHwFXupXRhPl3yO31W15c/m51J/jYlQcvtNcwoZ++4N
huS35obfIvpkttYvgDSd7nXBmLyXGqL3T8v4L+gklu+nFcmu5terGnoxVXKQeErZC543qJuF3Vqe
wzv/pc/WJBzmIBJYq5Cw25z6yvFE8ZtS7WoE3IjB1DwLHuuIX/BUPf2FhacoC5dlz/5IAZobbntg
0FHiw6XY6W7y1jYmCcuq/dEWNAMKkEAojp9cvyttQyFrabfiOF/OrApbYB3EFgsu8SYQ7OKORdwe
qh3gM8UFGYAV7nytS1SUAakfBypB1Vhh6AyvCCUYEVJHViLfwXQVwAdXcVXuTWd4KDw3HSab9YZN
L1cAJiUZ7nlRNFnGUZzQtf4QfkCIYaLbxbHCKRUNmjxEdt8pMFZX1dnKKp5ZzLaSGVvsuIVVRg/3
tc6FGk/OOBo2oMpbkKZgqcPzwS5Uf8ZUWEAXJ121Cleiuh5mnLGA9io3ACP0LaT9Dc7lQLEMFYiv
AmDFxq0ee0GmAfsVeNYLcSNMAfyf89CQlQKOdQCnQVXQGbNnqOkWfX+2/taaXKW9YT7H7Zh3wwxB
a43tlXUpidFq0hRF4ac4vt/jvxBQIW5Rbqqu5x6+RYtUa1FTbkvPtSrIsqK4LgDPBB2lewkfdVwa
8/5svbqnhpRPwEomDjLetnGbsCINyhdOCWjIBG2Tz5m5LRB4R2Ejso6YcHSIZl0hEaAR/OnmgkYn
Soc1dHBdWeWZtS5QHdHAOXOyd7qsI5PTlEANtO0/XH0VqzFkZRaJ9Sxzt/7jmOIB+qDEBFrqh9Gn
rko1mzhGuvQ4yAHfcASO/pUuuwklchHLiJ0saNiDnZduIYg44oye/Q0h+n8GLB6X9RskT/XWWleR
AdYfAU64piCZrponFCRVy8jE4aXHzljvyo0Lpep0phJgaZTO5MSCKLb0ATbnLTY+rZtf2FCFfiyw
Zv+4HtYsZ8OqoRVMQMsDM7TORUJpJiaSLfmT9TVzAfkdqR0Ssl//xq6KsKrVXl/IGtEGLOIx4Pos
bzgOkNJkR94Fu4NDXXb6WvId/Q7J21OFRDXz3BAZPNLzU2W0IpFocU31oeSlgiMHpikASSeH6vJQ
OPM3NZ14E/EYiefPUe6vrdNjhAKC9A0GVtLFxpxZdFYKoEzNrJ8mIf3kLuh2ryWH3uNZ6rwkyMLL
7226jpzWTodMEf8rzOBk/RvkbIeOQuLWS408QPVa+ZpVvf10M/H0jLh+0m9uBqoYxgrwuxN3Kotu
CoVDRnrEL+8/MQUH4qhvH6m0yle/uGxbIIjkwb4UfwUO09iP3fKk4VmZXxMRLKwuCAVo4KHtp4Lp
mPtWgoAnI8dlbiOP4+kXfBAEwXxIuJljb4Jg50mDpESskVKGPz3B/Trp+I8mq7AP/dNQnUlqdH+J
c6U88TAwxymljps6FYl3DGvtvoCG5u21eA/fPB09u8UGKn0D2Q2E2TAbgThXRYYeRN34DpvemXGk
oiA4DAGo05pf4lpZ24+jZVaJqmpxKRfDzX48jp0WdhCvV6sNExthaGKBA0NlQJaM94G0+PZXwv3e
sUMXykdfbt+nNaC6AN9WzKwqKY5oZZT3rF5RoYqWPVOkWF+6+QStp3zjC7G5q/QOU4jUITnAHjYm
KIbDb6gtPIY3szBn+fKWQhUPdXvylenenu1xDr/CAVkKndrPGuNh+quIA2OjmRYovNsYZQkrhGA0
SyJGbUlkI3UC83WLTSE00wriqCY4CePdbOs7aJrUGwLXok9SmAQn74WrPwoBM5Pa4VCZhEkpUY/t
y1FrXg4paRwoZs1GsaZ4zMSTqGtFeJOiSsHwskcwhU6PLcyoDB/D2BPfvOjEURJVFlsKU7Rs3rQF
aKa86D6XxpvhIkyw9lh05buZqT0XFl4ysye/iCcRDtEqTJUGUWQ6fIRIDlpOr+67QEwO52VM9Tvr
zq1KLkfTrinlOKsNJ9ZWFntXdPd81WDQ/3dZhJ+H98bPWEh0ROVqR2YZlZOsn4aWXT2p9Wc3VSF2
v1A8WbPEvj5II3VfNBIrHTp3ve0th91fobxi2P3nJF/o5y0dmaQn3lFx2ItOzx/to+eVp+ynysTI
1qOSM+il2NPeKYPiveP420U4xm8v/8aY37KgDPh8D2Ag/c0WMxPHbuS1nvQwwlfqpMtkWGF7aNYd
9tgT9R5sDzEKrUF5N0A2PgO2ksV73dQCWsgpJ+uT+gN7O2MkDditElat2ZU8N9IhOOpAQdK4hQYY
MKrmZzHv/KzF+5G7+9JYPQEiqLlk/NOGqMshjHs3Ma8tgaZv1+QhPb//5jB6g+mUjE3IeHMtJWT7
kUAUrEsQMEtgoXVVeAvR0a075vZCSR7ZyUu8g49HVH97wSiZH88e72BMhGD4TZo9d9EkcnYTYeXx
dInB3/biK/MhPpOt2cy/U2qRE75IeBGSJqYrm451nyMguynOtnRq+13leacl3uGD1/OlQQvF5h5t
NjeQEkFhjdsyKF1qzA9lMaXtBxz+6NL9/fUvlZqj/MeZ/dGUb1/FZokIFfWp0Z2BWmVjd9GkY6n8
vnI7L3AdzwnmFk6nEuooq45cD0s83P5H+hrak9inqJeAk/g4v0hgEwimb0Uuqq004BsezJ22KvrX
jdsQAM+igdnwWcIjoweb4PcS5emz769NVIt1Xn5e3XDV18FQHG/nrjAqiP8jgmK6LXHRxJot7z/5
w0bJY2O9bjlJjsyuGazrR4ZChE7gLIO74KpCwFsQl83NKTibHVMUCXrk0VLmt13c/xhacRf82A/Q
nDY0Xwc7ifOmgl+vvBGXfHavE3OWPKPU4zmHjA/p1BT8RTrsHOO6tS/QIgQsboONUoBVgde2gnFn
2PXHj51kwHHDglxIn3OGdefkSmbBDUQA4kk+nVzgzzw2p5NoY/Kqv8I9QCHTsPUmacKNDtoTFPgs
fQhoQsY8Y6GZ4ssQlS9Y8hxS33ems2R1K+V9DWFK0v0rpqlKO5nqBJOm6sRxW3lv84QbFrKz2dtY
FzG0rD1TosTXGSR2hvCEAB7BpfUDQ2kOlcBYWRS5n0wiFIDnq8rv0ULbo/3wW27+LHBkQNcYHoex
/lNNj8eJAcGRPIrNeJM38r1avn7Ix0D9K7mVefg0Xw/NoxmlGSUAhrR6DAu1Xdcuw6KwnMZJXYdC
xvP4CTNtVswhx8mKtDKKrvgENQxVZ4u7F3OE9XeNqrL5woF0vetXKwk2QJv7NV3qnOGSLusyWXSi
jyU405fd2/drYW+Q9p4Al7Og2mRrsStYalmBvRTKKS4gzpwUCcKnCUL77vwE+asC/sxAfH33gAH+
iVnOa3hhO5xCmCCE3dh3GxIjvZS2bmRv5N2/eSOhxv6bj3NYjbG76duWiTOyQVnl1wtB9VgnJCys
1EGUHAsSRfzeYz4GagVN+pyVhe8368QN5pBUhVVVsU7uriq0QuVKx4k2dGvbuMZxCzZ0u7Ev8CWJ
K2SPWa/JhgGFJfyiYJlnELEWAoBBJEFhmJnbec/XkuqSge0e+G0BneGfKLB1wPpB0MlBVrtuJW+a
FhsTr6MkGP3BggS4+Z3fKr7Ld0P0bwX/0pqJswOfw2ZBQaWwAZrERXugNVRwAfTDngsJWafRbYoH
RsJWQnwazSCuafO83jT84Hv7ma4v2tvaCpyafvUBto+2q/9lhnZwwVIPXmvFdaobWWB+HJLJ/LTL
AKMzv44qCLrdSuGV/i/Ggw6vaVbtsqs7HMVCrS/o79NrGh+xuBdVbD7+vGI7ko4icJcpg2krPWJ/
lOl/0Zu6RiEvPPQ0VzsBwq8AgZQFYVzANpbzATPZ5zlQYgdnkJD76AiSB3w5fBuLXOjb4NlH5M39
LBeXKVKYFItZyEnlWFY7BtUSR2YOzbshdj5l/9opP+dcKM0Ke+El3GQMCw1h/hFbr0cMrNPeyPMW
75MMZg3G4+l5sxTH9qc2PkvtpR0sXsZc/OqSl3AtsVilDmB+0GxsIREeQeHBrNjJ8aZ36SgpC5sP
AZ4tbE3NIbpUvbX2+UM9fa0S98UZQSpKCwr38A21LYUQXUEmYA7FmsJGn1zydYTcVsCQ3ztN2NP9
zwyaJy5amLSmd0+g5AvVOoZfUxCpA3iz6Hp1POwcJJTRp3pYZdepLOh8Bu33s8h557zEn0bOadxs
QZXn7vfiL3AflhvMNIsKGO/CAhoLwV5YIkMm0nUtxAFdc34wP3SdnSzn16FKZP1XSBdwLKH9SL3q
F2nKaa4/qhSNUwlWEF8+ul6ruKD90cJj+ZwdYmkaMNUelclEGgYFqjEscK2bsn2sKU/EriLYzSxO
NJOJG5y8Oqy+S3H0/fGq9bTm/Je6TvqUjE/yOqzY6ua+CjCs+2NXE5Q6+Zx1cCaSZmbu68hk8oBn
VpQ+xWx/1M/c/4W8qcPqo7bCg/Lz22Gg8KlYSAecDrjnDiLNruXM/wLVXHj+k6iOm9Ghm92xvKq4
6VtiNgvfyXornFLpzoXPg5tIAMXcfKgLpyBBpSupVnBSyUU/B85Tpqqswwtu98MoM8clqZoh2ywi
gMlRTQ5/rYMq5WhlEGp8gDSEIk6jO5rchGDgHRUKE9zxwTlH3Y9Tkr3PNeQzc9NG1BhBqjpSWXuv
WoqWuEM3s0XhbgsTEi0YoI4DdrAoCj8uJDJVvZ4BETG6qXHg2DVsItHCGHgVJlc06lqAAxIKrEfZ
aX9aXGV6DhtJBOYzPT8yDphasFj9OCd6bNlvv8NFdA+QKFkUpyBPsyzilaOI+o3xGuuzFasaalaG
+JYqnp+4z4ltT2SpMH7ywUGLCE/OoD7Pj+FhMT8Girb0FCeHWxdyKWDaq1f1d4fizOwfYro/EJNj
dPMRIF2QHmOAyxDkp9ge/ocb5D+27nIlh50HF2GNPNbLNnDacu/DwswlpYGor52+ZNBUyUhcnRuA
2cif4QI+WX4MnAX1kpyLUUhhfWkRPnAttXU9woUKgEwn8lkhfDx4WpEmrJX7RviwGzi0qTINieSx
R3VjOEwDZkyKn9BN4+1kcTKNdckfWH3iihcJVFkMtrsg3EoXiqqXlz07PzubuFOioqK0dNIYWYwy
oq2veTfNmLfcWvXs/ZRKh/3nNZil1et5aryZWjzEjmMugMBthQfScuL3T96Eedezha7nY00VMUr0
Fd6vJ/DBb8fZUVKKcX6sKE3uR10u6iVa43JLtpGCXukWISQRO2RbI9bIaVmzvt0vxGMr1OTjyzTZ
esKzycxxCvvz8uTahJkKbZvHt5c5zo6S6NfABAh+ZseQRrZv/vsoi/MhOkFkX188ZHyrqEOjVWA5
b2dhZIo5eLGNRJljkjl4/lhkJlSON13uaViDzQOJPs4zypskXhUv0ZcqH2qTKJqV1eE/lUVjyc+K
Rxoe3eKhI5v/OPNOhwX+X4VW8ZdptlimrjGNyVWxQHY4jpusseJt6R46U6cLFA3/qMaqZ4OAPLrk
KrY+71ypAgPDafvF+g1NYBKu5VZCV6tPl6pdfm/aPflL0RSJuiIFvuS/kv9tqUtSLBqRu2YboHYf
fvriTEoAKmd9pxLTbmrV7S+omKFJevgSq0/F4Y+I4UysKCkTcy7WaKfOszz6cgLwYSSQAXC03K5O
OeTDXHCj4A+QIAzV1aF8PWAErAaGv8a9US7Yj5zEvzYBzttK+EZCueBxY8TwYu9gCTVoTt2v7SwG
9MXoX0NPyADRZNnbsoqzlxiu9tnS+DjmmqDpri2noRh/KGrxiaeyRcjK2BDmVbVyIJbthU0f6JsR
9voAdHVoV9EF+EU8P2R8wqykzLR+BR1e6DKl4e5rJTG8w6mZ0NeS5furbImEv/2HX2V5I3RGktGY
Lh4Ciq5+cl/8QFofuJZ4ZABHFFG7THnWdBOdd+DmA5F86qStrsarrhPZcg2BEg4sJghxirhv2/a6
nHpRDISF4WtQOhrlRW2ZZ5pVd8g2osvgptpbN2r+z2TM6YzqEcLrBiQFTOqOh+RtStSlYgt5C/WT
RidNirXeJNhd+R10DhrB3TYP0cNLtSjO5SS6UMrQnPmUZhULdanwt+SWsl94xGn/6XOlJSGv4cqY
M5hMOF+v9ddcd0mj0XKeeOoQCBbIknavjmvHa2OWqPPhieXCaZ3nnd9kzsEYfPf7w8bccofkTouN
YxFM3GBpdgwW5OIRcDxluahsLTDqvZiCkFHsfz7OuJOILnbhibFUSk0AQubO6H4pNb7lM+kh9nhE
QTEW+bSYd1kPwR6+bRwHj0hCOiLvJQPM3/C5YqfhPZ4Vziu2N17Pf1Y6q3xsSj5ddrxSTtwiKcBe
3Dhfxuz/4jklZfk9+h4byOp+cxZR0VJiKExshPUpgNP1qtxA2DcNx3WUSCcadoIhQnsiHeahlzYu
vrC6xxxnd0nILjyImvmXX0AhhznuhrFyJRf89dD9aM2hrvtp62TmwEspJuGQ0lJAXjHb6vHuzYmy
aqXez94vuBoSEKgH4/qMcHYH3lOqIHmeo7Z+w1e755CY2KL07zPfp9Hm2zo1oCSXzMkux+wvkUXi
IT6wFvPwtwa7oZYP1A2tuTuCyWE5NceIpcCHpZdKazuNVlLlpjH8Xe9uTZQMYrcARgiHOF6oX0KS
2LfB62h8verk2TFQmpF5rKkoBYO1A70pa99UnpUJJjxpWOJf2k2OCRuNhq6URqXUmcoP3qHqyrrw
nwLNJoEXSB4FVrH53vs86DDsxJ+nhD3y+EJSdpUCGRBtRM0K9AxbSVZLBXzYBcF7nx0oKZI6ud7p
0OjgerOt9EJA1sUa8MAkid/qORMb1ZN3QdF4WvMqhlMdizlmy2Ct/cU3OrmBDG4HTHxK/vSWYKa4
Y7IyCWL6Kd2J3YUZF3ws7siELE50Wks7We2wts85uVIewDnZTAw496W2kcLxdla16qK14HwEOI0F
RH9UCa433WFsStuhiVuHnRPgCzltSMOwEFgkUJZVnHcJqWkXAf1j9Rj/oYe4i8rFaBPkhaKOogPZ
pfo1JsOiOTQ6lFLGO+dBA8AHCt6ncsUOl8g+NFB5qDrXhzWiVYdDeQVNqU2IkljjVHYJ7g/RBCZe
uYYFhMZVTOaenQrCmlmpkYJu0uJrIzjm8ihFWERThwC7WQlROkQoHDgjlMrp2IpiQN7b91heUuOO
YYhAT5z8Nt9bJBu+bejWL+1a2CCd995ZztsXe1uf3qieg3fKFKKA+4/WOhDtplFWKwb3gGaN4JPp
SLImIxGNb13wm5U+zmVZjWJzy1+qLYGcDGbLbqvStjfKC//D6feNclwL9gVLgSxQ7OPj4a9dUyI+
oYNpR54DYHTkqs8hrm47CaASRIM75S8WlxiF6IQOTq15FUnp+C4p/gYiR+inCofPRe6nxKjv/FYc
OyagXFzU2TvQJJ/6kDjEbfAmbXwjwu0pLz6dzP8Lx9jp8jNm4Y53YMWHuV7D1HlyWOerRCYmxh9I
LddKQ4mDRDvVqDGnRBC8uXzBxKdYjM5uZBlLu7UU1y6Pb+WKrpNF6H6Alik7GyZFcpLol2JB8XXX
vfoZsdbOzjBuZJ/5kcykp0xaP3/D1xxykdZqxs7SqafQ0K6TTaNhtfhSJ0G47dJ+5qrM5++Ix/r/
349p5gFmxFSWAC3yFjtNbOaQIi69vfr/3RttkXPvVYy0NvhYdmnv2H8sfpyWka8Bg29PwBXnUHzU
PQi0APIhpkhEe9Iuf1fF1m8SrMk/TrovV0C/x+OehMFLWQk77wkJp5mFG8i5mcOG8J9Sf8ocdTlv
dQDAXxYDp7rkHtBWC98bFSKUzCXK0Cpn1qp9B32RJOu6oOkSyrvOo/VlFRsy31HdpRJ/mzdt4Ibz
4iGzYAljQ1R03Ls2q5hU/aOyQpoKAkLJXNglCc4qlZXVSVeGShI8UdzhihS9rL6rtopdB33PWAsB
CVQuy83PAgUHvHA/RWCcq4VPoIQHQAjuDvFL5Naq7PiJYEB2OZu+fJtpH7ZYorWP5a2/blCaVoMJ
E+Ru4tyXrMSSyka+dfFdpw+yo13tMymKv1aLmHgcS0BK6oxqIoRGwAE4UjbIw+ihrV/+H96vHT5I
DQcros8118oibuPu9c0YKcsXjjwwSSnKV4wvcgvVnSCBlBdbWRolVs7cGauoqKNKSLs9JasrS1TA
DRvZv2RlefyqIDMiPzcVlvOrFBWDYyuPeWcj1zzcrvA7W18jn6aT4Iox7/kdayS9CieaYe7qwZ3h
5u0/GIaH5rw3lz1SkHhzuBU/6C2YBoPP+qngPiHmKmHkgKEWvC7+4I/9bnZpYRzkqiKDqbaEx9rs
uMQNQBz3BlKtZxtNtoY+PGdpg5vsy8dh4fs663LLLVFwtyAj2Wj9H5uIZxCmxs81jX0XxFvRjCxK
jb1mFvqFTafRf0M7vkLZXMV7PB54C4wrviLbDOh34PwHSe+lXPEkNEdPLdkncvxPCUxwx5wTIa2d
McAq8Jng1yGBlHR1VB7sD5XTH9nNmN3QJ9RLhqctiRnZv7C8ENW+KzFgcS0jazyOyttcM1PeXS6c
zOmlo4dibSxIvlElR53MPAwwLpSxQ3RTweCSMnnb1kJpRl+XXdsVN2BGYY78s/dwBI/cODzc2HAM
gv99HDKerTmrFXpE56+7/CyNArlaCcos7VEFhSkFT5QgWx+UOY3ZhwnbEUcWqGzF0EeHI+wyf4+L
WBYCEL9gscQbpSOZ2cZiPHJ9q8jfOcYyknxsOxNwArj53Gv6DydGVDHGVUOWsBmR1EOvnQsoC0MQ
vQ94s+NVf1h9ECufQY8l4Wop2v0Pa6afh3eUM6GHfGQyu9WPpmNmNELXqvWI0zdzxKuPznTYgNI9
JwNsONM/h/tGx9Bu2C/IgJZA/RDphyK/3DJ40M/EYxBYP3wicSbuiRTaZnK/mbqoc+VwFaXHS1rH
Zr9w1FhSlxd+fYus1ngZJI+fzqxweo72DEXWOZD+TUS5QDXrDlyde0S2csZYHxSfTIe8LEq5UvUB
oOMNUfZ/Chr+H1GVCf7/vBDslgBKuJgKgwV/moHSIyEZvJY/WSVfp+ReqF/v/khi+ihRTnE3CjOh
QYCtS+ffRAYAIBGYgtcdrGw5dhsH1412QOeIDeavU0eP29vL3yijF3mcCqPUr2QZldC0S0eY7koN
Sx+5d1dBdaVdHZq9Eaez3LdKZaZquWjIoA6Xmn8XH8Zo2WT3KXa4JQPOW6wFvSWXz0FS+DdbW1nC
RkvL+1SgU/kjfZ9FHea3t0SlvmPmBonRq5E31MDCLGc4QYZA+9dXmHJWSGyXcP/n9xeCzfyrqFvX
s2hnhtA0mggQRaVKA58dtTOBICDebEAwh9BuUyAQpTuOwhL68Yq/BOJC3YxRz88XkDHchxUJGYNg
x5kK831VaNOLEyl3ozVs/IvCU7En7qVTStEYiCZEecG7Xf8l3Q1h4kr8hDwTWlxNfSMRmiBKJpPV
H63UBE8FMKtN8+KG1X/NGLHe+4ASqc0/fjST4fREyusVQ9lb6CS4pkoYzAwHWEacdQZSCISyeyct
k15WG4oEeaKj1h8g7kbSYgVueP/g4dHpVC12Ff0gzzxICN9ABQnRZ9PeMMWvnF/NcFkXSegUlC7+
XmQr7ml1kUDh+v2QrWsNWl9l7jrpd0RLUJx8jOBaWy1XctClV6FGGM3dsL9z6XE3BYdg7isBHS9q
fPbFfnjVwN/tbnpRoCr1RtzR3jy0BHWZE4dg+lXYm2T5W5hPoyH8lEomcQumLVduu/TS8TTWiWHv
0XLuSeTHfUrYK7wSPz7bl0VhKqb6Lv+QQjoIm0LDIB7kDyflC6fGGaE5dRvHqemAIU13HnXc9Vm3
VwKz4nAyvOhh5FXsiRxp1Xf/oKU6/AwICYsbPUUch+iO351oAMqtlw7kn0SWkaNeS7a74/JEpvU0
XvrYjr+c0pslZLkPQlWDWkpCLqheQqoNvNNw/ffIkpqU+EDS8vnoBDD2LvZR9l3013/87lz+b6ER
N9IhtyXDln7yGyljwTiKnfJkywB1aspzKFIWY6FI49Loxrz1V38g0Ahp7lgMMfmvR+XH+F9uV6LC
+WGfcreoEU/4UjBvjIdlC7rvEl/8+kZeLF5ZDM53z1iYYoyFrnd5hgaCcCkNZSDyRNXCsRPgI/JZ
p1gI5YYpQNZ7IU5JYqlZaTAAaWAcZWbsduEfLzDFXuwORQn/xRcItNcdo/ZEZCXHqnLL95OEsg5K
xoHYECSTMr/Ndq5VJdp1aeq93E+IBgpBp92+n1QYu8IRGFKQtO1Q6x0PF8D1dPF4kT/yDGcTdKyR
IcjtM4gIUIMJhkN2PotfoVTqHuhiLVereKU+yngBTEs827G3RYYUq/0k+DxzdsCeVOfMRjb2esJB
791Uf3mtuuQHlOiCEefEqxkyMVUEVdT+USRrXvIYXzOVG45MGANbzKb/grVpMXzqEeQWHozGMZUS
Qvtd2cmjdk6qiHdMuH+zhDMqq23qvvXacNd17PoZUDCgqxG6GAVFHU3q0JH3aw+7FsjEq3VPsnBw
FhF6F60rgboROLJ/RjUTsScqzdJLdSpX5SkfreGrelAWNf5aNYNUYCpIJhgjbjkw+T+ob7oOzoNo
HC3IdubEVTq30BxcL5rf6Ing1YkkMuTMJyVPWPEkHnHLEo69Wr9TigfcIXuMukGZQ5fJ0e7k/yHo
gcpJD6ULsKHtLw9QM47fn96FMBvb2X7Hsz7n7+9c8TXw8XqXscKmTDSq/kccQeUMtX984NzsXtEW
rBgqd648QMORSN1EUPTF+rI73MCKx4xD2L0Z2ixHxYCsVZ5xnFjI8YlnDYZSuMYrRTq8WGlavFGW
hxemyoL81ZLuaw4nMLwTJCQqxM6m92g4MKBVNzSGN7nyvub3uzSxTekS9dEHxLqLRVG1TunFnZs4
pl75ikh3sRspbvtgQIejWhUzV7kfjbf0aedeBJ6QWU6xyqIq5/z74Qmme1zuvxNXCaYbGAumdFVS
NRUvd5Q4GYWe2TVmQILVCDwIz89Zoj6xe7Hy12Ml3HiFfAZTGlgxCX+SEE+d0VKMgdLq0Q3mjOru
jO0mt6nh7h04Yt2e8kRT1B7ijBpMQ3KVFnDjpdqS06EzeWn2EXvvJ3R17xPurG7CGBKYkjQD9O/y
TGmnEPLPouJGUOLQWu071QdAuxOjPNZFhRKBNs/zW/XJDsZcMzEq2uwOTdEoVDRqT1cYGZNtVVUG
+EmIqmpToUdTV6dPZLfsqw6sHBUZsIkdVDeTbDX+8pZHA2lmxReinLfnp5RYhz3UEAzzQti3PzMv
tQctHk20QhXSrnOSsetgD33TC1zXDzakyijKz6LizfjveN1n3eJPcKNXn0A+r7X67j19eioEwQnd
XahevRMEdTYQUodhGFPQq/DkFl52KKpme7IcBqKM7+ER2Lcp6NpX/fmiQN24LiMcssX4eqSMeYRM
EfonkUfSx8MhqRNLW7JLW58gbmlN5DoYdrGBlalkQzkzNcI40nLYRzGQcWJ/GFXyaFuoL0P0jp8b
iaXtM+5AVxOYZAmXw6do7NUVVeqdxMrOVDmEhtwNQV9ZDQvo4XLxCBvmEaBMsay7Kz1Z1IoQu++d
Hy1ao/AIAEFtB/Wzk2b+KXp/PMVhS1FSuYIbZKs3kQqNSatiNu/c3j26Baf1oX3zaqzXpod7ae1E
AkpYRpSJo/6Cg1hsEGTNbQ32nSrUpFvFX59whEG6RKWcLvTB/OzPTQrl745oc7g6fsUTman1xt48
tduHki9CVpX7Ex18LZznNffTCaWohPTQr3ldo+onL8hqBi4Bo1FHP+rFNzk1COx4ogsCSu3EgXIP
Ahh4a7akzdcom7LxXNOV9vpDRsDfzsUbSokrQJ2rEM3hb1Vlsiot+pHNgrD16HitQxPGO9gcNyx1
pLktCeiuZF3IlE8EagiPwPq6fnhZF1UeDq9261BXcjuvPBa4eZ4B9bkEVWb4No7Hd+lIA0G3ej4l
3R6J+efU6pah37KrIOY63kxErjgUMuggUyLYWod66MGCAiGK7Hao3mMCbmkbhb7yCN52VOkHuQuX
RIIGEKdjCn2nRly9pY0O+QMaLdSgyeivE+yXetUfGF7pcfEC05KRCTOzjFjL4sazfrf1izUim9hR
rq6IOAUln+VlLzH0SLkznv3PIZm5nIexNs0he3HguvYIx17BYqYfEpZjO7sP5z2wBHP0n24vtG4A
5CkNywKvvfJYpfyLueWTjzg7oPrDBBHn4LVnwKB+qHjsTkJQ7gjCl4WeGoFOQUU42prbuujWWwp/
8klXTOPc3Ss9CYLPy8pnMVz4XEWkHLZ6ib+5hExRPp/MshlgEmnnCjFYZLWPQZxCZEpnTQkZ7UGn
rkAP2AXXo1SXctwGYmlRLalAnz/RhH/HHMBpWKfmcBaAfg8mbbdrHCcP73OJnyQtDv8qdDl4lpJh
+mQ6VGimgl1Xpu/jxZA8ek9FcxUKIn2MgcR7ouADCVixEkHVeRvuTY2hw3ZV1eW0L+FsoWmgaoiY
41ONgmsUPCD3hnS9i5CVc8BekPENfHMROcpHekvV3+XFKaNle9kJ00OjdiCv7vt/HdWqktTGNlWx
TE2Ox9uSPdS0nDX1T86Sj4fURCD8a/gyUWZY6+0jAz7k8iauIMPa6fzK/xDA/FudnHTREQRZr+1U
h9tOFDlrbqffQkUGXwxP7fGSDd/OcaiAu5UA3uymhOpYQD6N4Qf/hfNjwZ+vvo12My04r3RRGdar
Cwf4uBCzoNj43CtrYGM4oUvV4slMYnUuHfguWX7wQ9HTqMOrEznpR69Eh09SNY9Yi5OEftIdRotI
Fp+s5Dyn65K07vfB0vRO1fYCsESZiy94ERoUGkw1MCq0tiFPnCFkjAt+90evN+UiiOybcRDlGx8/
jtw/bkSupcYKK6pwAZw3qtbqhFopo3KhUo343DpD/AXW5OGZRx/+MdmfJDst36f5uR3exq4tALDq
EwxeXDJMiOfRVjYDwiAdhyFEJ1jD5538NLk4wwVn4xtjCYXWe1Ql0B4acQq32LAr/xCcMmd/6zPw
gOjPheJYwGRawg/pHdmPInhLJms3cxPHwscLxx/xefn8iYMbW+wrjYE3OJ5mj1Osb4zfMeaxzd/O
CeVAkhFIv5L4VVajvfVaGFgkl01ZGfE/qNVBPiYWbi6l+6+TVDZCLKMlYAFv5jBA6yt6Ea5xbPn4
g6fpn0XUXAAnkSvYj7Ehbapc+D5FJwJzczts+itad6KnvBSk5DJgzItLBTnJ68A5dERWZcW/yJxW
R5D1z+qnROooSWyf8a76yMxZvVMoxvCHyKc1XB9tVNoD1tfCMUFt9T+8xF/wt1YWhQEQdGwoURgX
Q+wYpZJsMX3S74QFJddi6HOGHbETy7zzTYq8QGnvQtsml/r1sPdFqwJxCmOvo+VQqmuI5UDABk8g
XQauYvAzlZr4cXRDRPMjhJ+qCLj+W+ogSAY1uucaVyykrcLbC2CuVYM6SX6SL1KOeryeZqz+AmQW
nzTNuCiXBQmxeDkHMh9Z1EFdt8g6ltFIjwsf3wtH6nTXn16OzFWmW1PPKp1pfeAoFQS7zSr3wgF7
TVpkCyY2Us408q/csM00ng/axBAuTPYHq5ugxUEYlVua+iBIgqB3TjGoRfYTa0fJdfuhd5Pw2Ne0
OCqpG8ek/dvIiSIv8h3lR++bZCPqZVKW9MN7BdE0H0HqTDGzXRl8SHDb7A2PFU98Mcsy9H7zks35
eR4xmV6/0IvieWnuElPpfAZYiAT3BfXnJlic2qpHisbMA5U8i0NoxHiGbQuRZFpjUscOh8+OWTYZ
ACETS8oAnmRFTCj0gBAr+ug0muH2y+mU3qXAsv7tq7bQOzJF9lGcFPGlPhxGBmBm7ir0GWlDjEZ6
O+SQTVGm3RGS3ZFAGzzCq3KPWqmRzN+DP23sFh3o0BdyJ3NOAugy+ST9pvoYYuvr7IBE2xgxxnJ2
REgkXnp+3hnjiJdwPLFCsh7Ldk6qe/hwsSzfTYov/14VLZW18U4aSWZ7wixl13ve+Q6zb6GWzyLZ
dZtRzPhLfaqR9MX5pJBDloK72hBYU/amF/yLT0tkGb3vs32fUqACaAL2ICGVaXFCFM9Kz4trqAcn
QlezjKagV+e3c6H/DhZjq7j8mfY6ZDXBCC3OAOuElW3mfp5le7xjmSPZ89z5Awo7fyKO+jXMmZUS
aBUuumAr9zko7FVe2GZARXiB1VrnAk1a0EJo6Srx/EHDSNSCeNMcrTnfdwzYw+5XJr4HDRkOnWqc
5ULNs3EN2zUu3VzIM7fI6gePzpsUDAQDDZjRGoJxq8/al6iBPcq5RT9YWyxLIil2PNVm2Hcz+5ve
2xZuAVVFqtNnQDb6LO7ORnA15MHaPvoNi6GhJaXsrMDdyofw2PErwNKCK9R8uazwuB6FjPVs2Mws
vaZqb7rSxbZzriCevhuQYEqWlrsZhybEFP8xGWnCqIKALbDAwqMLbwJEs6G1TSNJbQ5vVH090TOH
xUR8jr8+8VQKXEznu1HHEdCkem6xX7MdyAr1phqLzRgc2XzO8hjwTB2AWeHlLCAmHM35csEZHDSY
FMtBt1O/lNyoy1tN814XCbyQ3SbbFJQzPda6sQ0bcp6++pUnbuCCobmzClTl/jxHOIQRCC6WiHwi
0zgIQXt50DIphLmt9QqBWYPjXdncm7ycL/28/mDoDahU5EOX9PtYZLMCOwjTn1vu4TK2vGoQ1C/4
oq/WZeOs5uLnI1uw7s45f524Q72we7m264nIP3nzlikuWHSXIf9BA15/iq6WNiBrZoGN1px07EE7
p4nfmpU5tPGvlzgre5b+oh9ulQ0XtHXQF/1UPSivtJyuanGVGtu74pen07uC/uB9qrVxrJUJCeUX
Mjw1+wPu3V7W1L9ir7o9/bdHi+7dls+8+Q7Yas/weFXQG0Z937k6SzGGZhQJkCWzJLdgqFa9xmlx
gc3sw4Nkbz4pt7v9jBgQzRd/KGjA4UCCa+rAnIRukwmMxqQTT61DcPbb+UI/MmoBOciKJ/WQU1hw
GwTecfb3ZnuozNLDHwghDprYKk0Gng9kwkuca4VI6qckPbWWmedkZ0wpzLN7jrY6onQFD8Y2SXv6
i0VtPYCmTyAJ6/pLCOKuQRSHDW3ioBchEgzF+1I0U2ktBNElt8dafcN7gkUqmzSNN/4p+ATA6A5T
ZN0wSd+9U82CQri2pJweB5le2M2w9cfck5jlBlVv4H0QZwVbGWESK7Ujb/GzmICJZgqKvuHPnrNU
qX8naXp8VSYRFa9yNKNfvdwXVTlhOV6xyMCl1iOlaRWtVUE8wkc39f0pYTS4XEbUTVVsIErLmshj
He3kjmtpmYBO7s0tVo3N3oQNVKd9dxYGyT4tVjJAYQPXagRNQy3jj+sDYlvIU35/pgLKSF7oOxa/
jNdnQXDSSWuapgCI5eJP3FpvKDZWQzK0TQCbYz5JpV+RwsIa6PbDRy2oSUa4JZTfY+C+aeKudfI2
OQNzZWxhyngs++Y54yxfyTgqB5eD2b0lO2uRdKoz0k8aaSKc6sOegHmehl+ila8e3VNwJZz4Xbrj
PdWbkM3fopaZmqnnl1KABKmk/Vnq1MVUwwOhClidnNcweEYeUKTkeMZcTiNq0jeSy7tRAHZea3O/
7zgUZFuGrMevQGX4Y7p5FzrnAma002QDsPpJ65Hm1AnQYS0RO89c7Ovm3GJjrxxBkoIQ1jCx+oZ1
jTIv1DlNVITJ1KpsP36wJiiDj9f+uRz132TKguszPGGRoDUEKmyj3DAuwbjzs4kZ5URmxz0lQwJH
o3o38XS1AVThF+Mnudi7W3abEVTYlYEyzB2FDQJ8Mgn+eFFPgfwNsQ3rTSBp6M11hAYhiDyUaGzt
Fao6wuyg0fJci6f6lcTk1dWbkw4H/Wkyju5E0WtPETyAsGWr9AYHn5pKS+1Ouf0N1Ka2htZC5Utv
Ngk4qk78bzByrHZxlv8id7yTsGadGyk9VBlPBiNCqSCfIo3PHrvrMX6TYtSa0qBToJfogB3JfM/d
Am/d9Y09yCpo5HBfKy05S6yhNCWN/pkiY9oE4z9JE3No74a+s224YSPvf0Qe39picko1SvSmWDW2
AdaSIYoTEVd87qO1xvVuaPzdJvQynRCiefVmuZOgwk/2pUBNc89llA7CrfcK3lMH5+euoCvZOgYc
nO3NV4f3y9G6rtK3OjPLB0Zjj/6n0dD7l0i3WAjhiY/FnrIfx+yOd1pbUyRd6OKxqdcFdGgEyTLT
GSIVaJNhYNYxxB8DqLvZMtwUWhVO0PfwTrcJAJ6int+6Q1lv30/qR8bwuyGdDEQWa6n1sPB46HrY
dFQjbEzM7TUcN83dIlOzbWjiadv1FQiW164ZEo7UPy8JlNHlAHSJAG1xLvPYS5IuUQRuzR6Cboq0
VHls9lf4piFnbZBd7W6EoqVCp3MdEi1rAgdnrOjrjsQH4bqTMHxaXgNE/INn9eRVYLcO6rlAZop8
Czc5KlfSR0LdtRmMS4bOwqFNf102SCd2PNcS/5dyS1lRxfwV7s2VBhUnXEog3dWgU52oZgFb8BIr
k8EejxpVYEvDvlU78DP2FHBdmh/1hnPtqUIl6Sjy2u7wQafdiWEW9cM3IsVi2UUK3JPcSxj/cqj8
QqksciYf4DVCqe85REjNVWzYA7ai28yPc/TuPRdUUxn1aV66vdCooY33xM4esij0oXPXhrQrNLUt
JE2dYjCZrNTZ71Zmag0U/AlA6Dux3Rufqvs1/jREL8KK7MPFcbB+lPSSEriZt7hRznysOkp6+nSg
Omw9x0DxAz4ZxsES7yoqKMKKrR06ec07V/skYkqirFlZrqgv2DZcg6/1MHCI3ORwHXS91hMZ1a+L
oHNcgdUIem7QH4a+zigstz0RLNR5P92UzFV3RvUXu6AhYBVI7hboq5UewH2VKsa51l8E9pZFm1id
2FE8GRk32utUwyDDQguFUzgRJZKkvoplJoGTdDwkDtIsQOX89B9k8P4mNGRhuxAayUrKcKknaNag
wXgQ7RZszL1/bxqdIRqNBwg/WE6J5IZcbUoVFmAPpZydPpV4yvHeW/3/npmM1jBaIBFRHSzD5KjX
LX/jhLv+k+vZrv0eXA9lOO4fHpUAYSvOXcbx9ZD/CR4OBv7aZ8IFh5+nuOMZVQ1PnrrW7qIVSUPa
KK5lbKxOiTcu9vL/9H2HdL9OzVcuPMaRoHHbB4rnRlg7K8oCin2xssgcmt/A6IGQS7tL8VSUTtq0
wzNGIp7430a+IWrGInLV0CssOUk1/LAyJCaqLBqYQ6NaTdjgv3nyNGN/6lvQpOAmEFMa25wg9A9d
aL2AWg5Osf5qEo4x+2vKifT0g0Jgo3ex49CI09UPIdApAuc221yz5y0Sczrh7cVj559Y9PHJuugw
+rMkDX4wI4r5tLOpLUs/kt9UfsKRWJQCMfc18LNEXbroexWZD2feelQtTYlJ+8Owo2fl9ZU9sHJJ
qf4EHk0Wsenznb4oK2sMl89kohmyPMs5IoVQukh64FctU6qg1ZSqnt4dRdGoSVCWUCeY7ILJJQWM
RaoL8ciGlY/CXJzw91+pEUXZDl+Al0lGUnDG1Udoqudf58orKzvFFr9tRXY/CFGz1q3oU1rOoS/Y
FvcQWMNptnBx7jIjKVrUCzvhRK29p1tn09QR5Z029UhxNpF0dVDzVbxS9/BwNxh2XjQ3jKuLrrZ5
nCkzGL1hUFQEI+atXloGSP92z1WnrmTt2/thLBdwy2iEqiNMlaHAFIHJm+X9Wvi2UvXsjnou9asV
D8cku6Wv1vv/I25cbGPP+xKjKf6yPdnwtHKJ4LYFfSdiMMHhSrKCM9tPFhVMBjq21qhFzV9YBx6d
xjS+ZxMqq+lw+1cvy88bEeOuINlTpXD5LAHsK3YthxeIb+KVybYwdjO34aP9n1OX0kTViyIZ8Jnz
UK70V1lcfXrcJvaDwH0u/CLQ0E3MIip8KIYBJGslDBAINRmAoHAN7jmcg63R0+P/S58XLvwm33bT
WESJHzVhMX2dLOqMjZyXnG4yqTpqpAkOpZsFuSYAY9w365maFpv6pC4Jycru09k54irB6dZQxnhJ
+52U0VhCLPJXtCexCTlCobDH+5ylBAzQQJ2ACJP4sMZy5YFs4bZ6hr8TZnrBofw97Ij+uMJyOB7m
ZU99B7W8Nqalw+9LI2VsdXudUcR3kTTo6pFKxZ9WCeWrHGorSNvpBACnPoDr374+1NTBeOE/eSVW
1GgHTcpCoLPrwFSWWk/9OgbeWND7YETC3OQ/M7LPMc1E3SxAmIERr6JLuIeebdONU0YVtYbHpmsr
UpVzgMkcZP9TTQXciNdGyuF6iQPUyNYo4rZLuXguYzxPCgGlPAFUCggkYodLoh82DJfcwTt0fyWL
UmHnFwj17h6l75hycN3280EMb2c/KKOG5N1y+lsLR+ak1cH9/cqy8h8ORgsnZZQEzbLfqB8iRqbg
KtPl4rWqfbE3xgVvnZryjTnUko+XJ9C0O13ES4Hp6OfnJUdVUA2a3vB6795Bel+O5BcEhWG/Sw+D
WU8RvZnlXUlBHdurcGUh66MfsGmev+eJBbf1/xkgn9OoBOfah4XOijHJMBqc1CwpNRgAevoAqOLo
tbqGeYd7DlAfd5FOmj2YIe8mUc0DaqO7voACGaPIUG7q+Zo2896u1yu7OyAp9nEtCVwjo8GVxz09
++iynWM8OxNrx/94QNeuzxDI7R/DJVrIOJbtek8qrodJlVX2w7kDMMpT2FxZHM8WcG0esY5B8D0w
+EoLplqvBTvmezJHPiti0Wjw8SQafEg7xSTJYcOIZ59F3huNLmYRp/SWoJId6j2VYuqZiEFCjyOW
fz0ItI9mEvQFxRA4yZaqcb4RK/JJm8SoIQo14E0yhG9GHqVVOJc8KvnRfexvMqb0xYYAO+v8LifM
pO9TBQNh46IfbENrR4PY0SoSPRKbJ0Ts6QCWRWuCmE035jiPaOBwjvxyC4xDJnMk5bJDe9p+7awx
1Kizrs1STdyYp8sRW7WDxNS1BxMabmIY+k2xqR8bAw6iXZcFTj9ANgpgHhGMIBbMI3+QNFH6LoKm
lQD9U4nNj35bZcrZO/bnYtcX10ECUjxm0dK0aW2QbkK7Rg0Nk0ZKWiRwT4SgQsQ5SNhlwP5Fteqv
ePiuyQL0fSEdd3hnzrWjJ/eUwddlsqH1rgXdT/l7K/JBCAoJVjlwsTFcR6DH80ae3i/ojfGIh/ML
EpMaSydhiBlqOuVonA4//CdoVW8ZDAU1D9jg1WiwrVTBlY85Ym2bw3fLZmHlkojmNyEYOZcNdovv
tg2xSs7SMt6IjY/EW1IY6HM8rl80/82/Q1LNILBBIb3X4fi0J56jXvOtG5Klo2iK8iKfTfp7gcfA
jmsHIZ6HZO9SLEENgobdGIN+sMxyfWtnSv1lzlZNXLrM20xum9TS0mgldPZsMPgdNzmTYxSiHOys
nRsdLYZ2UtKvjrYV91gefHqAEqTeI7v2L+PqliON3ftyiACgqvXRIJL/UaxEJAs3ZJXok0neFMHI
lXOSVGzQmj7AtokjyZpnnklmt/9bCjITyAfzg5HKatzIlSfO3flaVUzzq31YV5EVNzln5M9ZAxVe
rtcmFU7KG4hquW9uz5rNdGYG62jFM/3JMKpuZH13m1l6Eoa0vR1OJxdYdamlpHHHGjNUf5WcYJMR
N2JwjYdFSEzXoRQkHrJoDZSC7Z4aE+0S0fNaiabpdaS1y+03rffos66R1+oT9p2pnYk06gDvA7Li
Ny+kHAlCYxBG3KSy+z1GfMXA+mlebc+8luLchnG4themcezjfhLUHa8LQfmXRIzKIagi/J20EH54
uaYPcVqc5dx7wrJqTmksX/Il0+4YqBYdRTkBDSIv3nLjCuVH3e5zvdUixUn28Et4lyx0Wpqvbfrw
RlfyPhVw7y/HkwjHdwrLQ7RwYOrUAS7duKany4VG8DjleuJ2vdCnAOjnQCznnlisXq/yEBf6RaT9
PfX1BQBnrjBbAoxgMim5/gnldp9sYJyGsXFN+bCgrT89Zdt9Bz/n0WQ7kq7ZMxJ8uF8sKSVIImah
8lCXGDVEdgkqp5iNzKgWhf9uHN3FdF4tLFjjftF6ild1GDlWHMsgOgKejhZCjUoNX0fidpBWNoDG
aumujdOmHvZJz09kyMJMoTza/xkO8KTSzs5mPh4mjbZdjuM1pmW/73tnL2utk/5bZsXaU+iL7jeK
Gs7rhfy7eeGyOeU0GUVdxiHUpOjthszYI8OYV0oogK+IP6+c4akMzUxSHgYxQhjtfIt5wQROJF/S
m3GY6AslSoXkONH/54L/wWanUtH391CZt+ZEMUbed13K/mt+RGvqd4+YFy1x7l2PNO8uwKKcuE44
V4fHlY7fV7xQvZwbr4B3g1NgrUNIoTCBFrrRP9efw6BqU8wT1a47FQ1oKQHCOCH/45V1sYTv7D1j
VdloabtZNDJHMTbb4yhhGF+LSlTBawwleshRfQKtJpAlB/bgXuAcDptL0e67ybNjm/vymgloqo0G
qXDmw3idD0l1IixPITnKMFqj8JMmQz6sCt+vOqFysZRy8PziJNnw4CEahJN2HCQ8vf8DxNcAI60P
SQH/GisNGzhlwoH8Un0ek4+pyNbAAjR3F1e3vuVvdMrABg3YbZYPeCQbzAPUERBBBiMW6HwL5giM
ybC8PUDzuV3kT96853PhML4nZwNSC4WkVTyGKaPjwcb+l8Dy1h+KfVmfHsDleyGTjog38x1WtL4A
oBZwffeGcZ68NWxRajRs0Ocqi9+OZemUdoHbnqXsNkD8Uzi5nYPrGYwh/0u5sHhuEzQYeOu5tZYM
ZirhKSXW47zJwOjZJPP6yuIofhNZh1zL0JsE8vqpIFkpxLSvNmmjX6U1fRIqMoZ8UwfRX4f+oqVK
F7JVr7RtXcVtwFiVOcI4F8Z1hl4FiRUG0y2ep9bxJ5niufl05UNwA99wR4bpia8vpB+LIXXPgmcr
D443GzGaufSduPAWBi6Iq+sMvr0slLpbRSHHE0id1BgaFTaxte+gUC5Y/xAYUEgaXm5A0EhGnMrc
j3qEuXBIuQDff/OWejZW2w3tOOFT0yoSFmwW0WL74pLIUj12232Xsk477rpXiNxj5f4b34ad0kqE
IWWqBtaFX+lmkkr05l3P2wbUJD+kk+WhAjdajb1k6kpFCXiIIli4O5fban+RlkVuoqASlMjVL9On
bs7N1Mh4mLje3C7tPxCuxehSH67WorqZvuKCmTRVwDllcBksHRNWMurH8NyqrHpHICNrq9762ipl
RbqJcQ8eOoJn2iMFPUMZtFKxlpHWsb0Rvvl/1Y8C7g6THUVL2Pu0IATiba9aYMU9BR9JnrFNcK+9
q93v/mCLZvROPyUYYpvPc+nDmGngjwFc+egbf6YvpS/1mHMxv1+je9IfLEy88iAebRW8kW7OKdmT
OAi398YeLqGIIQoTL5+pFmILY6NEO9VNYh7RbuCNqYHT7XWEX7M/o1Y0e33/R426hznijKtrEP50
SSANbCKZgh3RX3U5y8QnTIAo4MnXV8xHYUd/fQK3IyASIABNSG1dw/I1Ttd+yLrn0qeokzmYQwNo
k7bo3jy1Ltm01Q+h584PhOX2f+VJXScXsASQGLOMsZvAidqKUMb7YFrlGdteEA2c+VxvAQrTPlHT
NYmzdyJa4mUbvwvmnSThw3qhKapJI8J75WmSMuh9ZnEGL+DYIBhSLMVFVRLputORl5Y6pZc1cvkO
8IwOW8irue+s2PF+sHQcSsidXm7wneE7PflfU2m/dv3KxlQzyLSx+86CO2Kr5RVgoB4IuJ3OtWQ6
PzVv1ayt6WWApPTwdEQhIq+hnbM62ONhzhOOLl1dlt1xlO+FuImq6hmAUnmj0Kd7SzTz+oxOk1A1
J02a/+naPJ/PLfOXHqCZJubsdhGKk7MIvIpSrSjPKh79In5pfStQk1S53fUjufvrSi5hDF/RMCak
+tTRIgTaFcdUEnaXh9o8m8+DOJUDpf51obptgHlhxvwj3X/uKNKsI85lD37h5uClVh5xQFeQRzxh
oBYHK4hWLECWH5mfRbmzD82W5XfgWjwGTf6D9mIIhsWmirbYgIMql3aeTXObgJHTAjq21FrDbi8P
CzI706BqAHgeR9l/B56A/cAc7Kqlo51IKT1WaK+I6OQzpdOh5kdzWAcEJzQedy1ddL8KoHsd7E4s
W65K97Wpt3+9qngvgot+PWWg+zzs5jomu1N8/5nqOaHlOcS6gVnxIH14Ql/CXCaB753VZBa5+mvg
ej3wtkNOOuxXjJueJFsZENT8Gep5E2bAjE7isqtD4d0jWeHkJSrRDjqTf0KgSikNGHaB/h9SXkPU
G6r0rwcLkh07v87aOXI5DuBb761KsOmPQzXrrGYz2x7ba11No6YRGUa+gyIndxc4/CIwSgC05lFM
f9ZLNDsfxx9ZXMkUNmzRzf/d2TrdDm3L7V2BYZ8JT2QaB2fdj5B1auwGuqvA1OeIRCwtgNvwFuT7
a1+g8iBcsCfhVMi0FZQ0SahkonXwR8Cf8k0S+dmUOjGCax/9ToiJBMVFNP0NXzvytM8uBcaSmFLw
69O0kFgm9nmW4jVZOA/a+n+67j64ZiQdhbS6pHutML2QqpawH5K+GLRyy3ArsnqzQLFcQfVDdtAT
0dOBdJbxObsDJs34Z1qopQbk2arEFytHzzOhoC9An3kh1R+QS7dD6fGqt5hMcWpAp75oFEzNVMxp
lsdQE7jB3GSALKiYzdVgjPmYfg3axV4uyUE0BykA8EQi+S06Cx/0A7dZmehdi2a/Np3Zhdg0u+DF
FyxMj2gm5ioCUDZcq4+e7M4MEGViPUnHFACLUCSBS6OGpTsvp+Jk2l9YfODN95ITkbc3hdk3TiR2
XxDk0FebUcEFbSd3HlsrUR8Lz2ZKIL6YrjnoPoSzDjqJ7jGKVB06UEBQZMRSCkxV94PDLwIMoi5j
2lmpHJ7sIsQhooB56di+bqw4CfVE7ld8aVQcvgsoRWXxHluCY8/V1ca7P/++Hk5zfv/suy4Iu+Gh
REu6hLhX/GB7xEwWXfWj8qtQbtYAwa7rj3iadxl7kEBFRIT8UAuxgtiL4nVUHpUG2d8UEQRIYyQg
Panu9x91AVBzq4Y/B2I8xRa4wbGO0JoeHOrQaykB2rmto/cy1h9cXXHhtwHQxvPAGQsDjB1g8unp
55/OUqvbSDywmedLl8G9xtmApKpsQeoQirzjSHv8fx457QslsclIR933FokdfmWoey5v5BBuI2mN
K24efjipx7FHX7AE3J3lNPYCWq/lFdx7/j8Pa2eSZmKYiqjq+x7RnaHYyoHYrvWgqhmOyrWFoSVp
Sr5XRw3wwp3wXvlUBu4M+HbP8hpkQ4cSpFrbFd4sUysCyE/ii4GAbdarXHRjS8PzklpNQamvZL9S
sd/zLRhJ9kKUdfavVGTURtkGF3Izd3duyS8wv8QbGA6+z1+qu53S1sIPiaQkluVZiOsymp2gvVi7
yok3ID243+OQdf6jx00ke/a2CWJ9/PRjL2s7NB/TYAOOB6Bdx3Zk4WK5h9l3d2Pc6WjV6w2KtI5i
1gWW4FCbm7x712l931t1XwKmyUBC6ri0yFOPIlFu3vxuJk2hpSmThZ48YJGs5jIjCtTZQXXuMgg1
kKPn6FbwfWfBBsR3glugetpY3RVPnfTD6ZsJ4fpD8WBTqRJF3gA1j4UpMjgMHyXsz7svamvHuew2
J3Nhgt112X6/AhiSfgI3V2nJFGYKOatFJPb1DOYesfvxija3H8FfRB0Cx1n1J2Xe9PtA1a8QrbBd
2EUR4XGkdA4fHOcUEsqVfI+tncTKQCHWC1QqKuO9HFqDj4e0h6REqAa6kxgMAX8pdRg8a6CMV7Gd
uckpO29Wa/38AaqLcUQfQWOxrGyQoWBdcnx7Rc9xyORRBCTQTNV+9PFbdS6PXvMHXDwCLi15nUaj
xL+5O+s3pYfRtfjRXhmqbm5ASPBuFK9nmnVDDh1ctd5S3G/dGjK+ySu5ZK1a/6BXjyXFyQIxARF+
bn5KvM6OqavOof98OtLcDtLtN+yZphBJE96nZUbBUKZ3tKud2AZ/Fk+52l9kgilbs/RWwy6J5qqB
WLEfEuQOhgUUBfpQtObgeYx6mOgNHCyP714uMpvA8XL0lGK48+3vUs2qSjJAND4SZao9XWjqOTmd
sTNzYLFNdyV56BC92AteSBoOHtKs5oSXWQc3/hDmmn87VpSWdD9hHzfc6/WhZQAie5XV/CfgHqWV
iRGM32rrkaz75L3ihwLgrPym1S1tnGjD9nBjMG36sP9yvCb/GvHYr7uCyqfI8CBHc2UfL9sOFo1K
6zYJL6RH2MUJufka/04wPCOyoU2ead0M1v2qi7vBkmPCa7aD4ynu9EqEx0tUwDLg42ixlDpjOHNJ
2tlw6mCE7do9gRE3xUvsZ4MF1rD5uxe/g925jEftIqI/0u1tkZqAwcOEMrFp5qQ2IB4X74hyB7zi
TZfPtd9slL6Q5tw0uW/JNuESlXCW8swYQ2/fSpyaBOpKVw7qVnUYA7sxHCAA5SJbIZTNAdGVUy5C
b04sbWLyj/0ekVB8t/lE0k9RpHHthzXDEp0+pdzFbFP5nZ2j1iDgdlVyKUTpLg44rVSJ85WtKDqN
DdY928T25CLLD7k6Xa+QiHi+3Oiif6DgMYYFZME1Ys0mEIQmlfDNEtFkI2QJGnsTEMc5+ZWhuvIb
mlvJKCT0o9vLQDjrcBZk53HZdc8E818ZVvHoQnehBLCZlQFIJnHR+6NcOIZcXpcU6pXEwirVeuFS
UO3VbMfB5Eaz4X/SFKwAbiPcFX+qumJt1mIHk/kR4kQ1CDxpp4Nyl1lLXV0P35cAS6rRcwizWWSE
AlL8+oP9rvb9RHbSHKVa3IGTJnqiu1HyR5ghNRsYCN1skFPKeNo6cvw9IGviWNdSz7g5s3N+1RI/
Rhdh1c2KeHJuPoM5oo+IFlhTd/rAZZaLFF/Cj/ns2F1LRapObe6NPlMMilBKP/U8cW5IM94xnzBP
DknBju1tN7XPPkFukOLP63fB+FX+5VtkWTLqigzZuhU9IjfvAdo/q42sWW2qQ4xuZk0mCx0G4mMH
phsgj7LPBj0KdImnbKZg4wBt/SCmhOvY3MrHdxoL9l2sBYrC4Onk3WRG3Nv1cRaVMxdhZy102zD2
i+43NOh+Rs42I3KiABK3sbc4dkenOde6I80youlq+b4SdxVaoWmbmmGxEKVmRe1xpGXLM5F7Msit
+l6fngDKOxcc1K14yzIfKgMU8OO3Z0dlk+WiUFmV1ZAzXUtc3tmLbMpI0opz+kA1CPvB4nW0xN2U
xclxkm5kcwSDrcWUR4iNvD5+42/znrkVK4javdivYrxmor2xPJ/A/MWClBi4uHDzsTEp8PRRMkbg
lj8KdZshtoFGNY7sxsUCWutyTeV3FguBDiMFMVHzvWHCEks/eIPWN776XTopVeUyXCdmar7LNSH8
jJ7jye5+n5UMArqT7pfDoa4E7qwjyXFh32EKbJhvsDguEH34S6KmHx2K4n+lSqS095NBxd3cvMjx
hbU5hGCEjMN4iAreyXXZMGViDGT6vn/Ea6eBAfqQlpcxZ5NFf03KVJevM4mCTFdsOve+CtLp1RYg
yXArNszErJY4n0G0JwuwmIr3OrSiEs3irdNd2m/2f5G2LKlM4PYXlnX/orJGqltt1WSlI/RUXlnc
b5K5jqF1bXqek4n6yQKlPoGpOqvc01jE+4fubwFHbYtffCBlANhpSdmPK8PesMjqHzNclKT6085m
CNuj6ypTocNi13GmDv6bDh95gGTa7wkoHy34UYAJYDruc5NcSEEduIpgyZ7J/OKJeGsw7cnmYws0
hrvzKAbYM8d4JBhgwRx5F3ohMjvAPjcnPO7q2zIPpTuZDrKysVjEoZTYjGbVNsRiSsppVYn4TxLF
lkG1+u+cGjrZg9ihkofRfdRdGhNao+dn2N0AHcOXHnnrHRRnhTqJ2MCLrvuS8ymD9uDcFrfBpSrM
D+A4Cy4Pn02NcCyUAa1/HEJL7FCpjxXwEyYgiW444POVR0q1Z7+kqL5Fv0THV/SP4c5Ctqr8qOjW
FXeKcjvCPJTdoc0bj+tkRx9zKPniRbKENbRhmbuevJn/Vu1qSRQlRwctHdTw4VoWQxrM2siluDO7
iEYdCHJREprnwPgiBK8CAkuKsFmjy2LzxqHTpKzWr+BSFQTVyALttU8G4mKiWZ0zkOK/2Cb4PesB
OCe7oz+/XC+UYV+oJSbE/0RXwxNm9PKG10jk/di4QT6MAa+NCwV5aofVppJR6nkPKQ+z+5mg9TGl
alUJ9CaeKQTXrbnMNEuXAMdlghztGTnygPgRX+ZA8mZfA9l6zvWlaqtZROF0gNnEHRtOlgh3iIIQ
Y1698P5aKG1l408zhQh/MEQobxuV63ruGM5fLa1oafZ7o3cP2sgwcJT+DgQP+SwMBrtwfNGef18q
45kA1f112UdxaWwjElHR8KxFICGB/xkmiHtLn+diM9Fk3ApZkUp9PMJS7OfBMW3yBSvE0c8w+8r/
iiYLVtxAYnszK3/+TEnuIhMF1USO/kQhZ8AaZx+yKuyGOYUx/oSNpuP5qk5UvsIt6uAV+jazi4cS
HgDNp2eh1F3ZKwdfdZUBqAG+4P2KEhYlWaXLy2iOkiZLa0PntaaLL0hfhJhG1O0VPor+cQsstXZn
XYmGyz08pwvdHe7QiumeJY2jwlFJv/g7B6m3jK7ouldnEYoNPmMyBqSXDHymNiKZYku9ytb3eVfn
NRG4xpVqDH1DO2Hdjc+491tY4/i7/wmVkM8DVKwaFo5ZYskfZWAYtmh8/B5SF0bjRS0cDmjDrbF6
qHXJJ7buLHB49rm709DahavgXXVqtDenYWzSDr48dydegsaIU+DqPzhyDDIXe2bSGSDWIN+6ZorR
hlDkNi8bFC3VWRkpvofmds0AgqQ1YSaTTOFiCZE5KoxeLYkMO/El/pJCx67U9Lw971eTfwmPzfhz
gLTNryZHOshYMc9JrHxQrQU6jn5ZBE/H/xvhfz8O1bOWb1f8TIc8eQDG17aDBW0d3MhqZLcWRI42
BKJPBqiytzRImPAGIS/YJe20udwuDJMIaTfwbHZRxemdognYLRlVgRK9eEVlxSFjiMrI7zmK97J/
nleqmpiXNtP/oVZl/q6qyDHRhk8MXeOD4ry1r13t1+oXjbbt2JLZvrI+1abQI0VBMIo8qXitWYAa
/P6RP4/2kRAMWNwRZQLqyEUIOUYBW2y2TQtdPpZFCSm5MIpdEAOwVAW1Pf0ajbdBMr9i82OGCuF7
6fhDH0yp8cLingvxgfPM1q5DyjNCH69AaOuL9QLcnczUUxlaRiBWFYiuGPvwC3pY9kxzpJGOpve0
APefuWV/0DTVRmL0DCgRWdlrvj7Tffj9UpZUz++5kjyV3Muz/4YP9ZfuOuQS+JLoK4NfuQ3vxJbx
4HiEno6yE+3KJvr4JhOfsCd9s4yOsiGqJ8g/iSBm8+VvRdKG+6pXhu2WIP2nMtYS8OO7o94bbyEQ
1ZrnWIQv64x0g3kjJnmgKncjxwHhi7TxQne9f1nL9ubx2177eQugT8Y6KDMH0h8P0SBZX15oSG0s
wiNyzId0kht1VX7aXIW6EboFBxsNuZkrKLFTcwhFylUauuWqkwmLRHkR13ygP3tteI6LZDS8cPBc
eX6JTgAN9pCmHZBB5ccdAgKMnYlk24XgQAZ0j6kMtmohBEwmFrBo0d8IGYEJPud83puWozPy3MCc
aarhzM82b50RMWvrWfBrg13PUxZQMw4RnjVZUdk7F/+dk1aY0JldBLEM4O57/SqtWzxn/q+OjhZU
pccOgpqkowyGddviQCLLMYGI/gacBejfNb5wdFU0tGN39KZZVppjvA/nfvb6xnBQH6XiZLxbONZJ
zoPOx+DGkBoTkMyQ9G7/XYIizyG+6K75u84JhF1oi8LCPh1wwlWBq1tdcOW+J+zg7ab/o+BpMkRi
JtAqS0A3b3BxN7L59I0XRXU+y4yiqTEpk7cLpFlw0I0cV/0z2GapOSagFMrAHv5LP8H7xOhUGdo4
4xCo01qbH6vKNBEcE1LJU84cd88J0xZvvKz/ZbP7a6+uuRsvwbC3sj0Tax0CvUgX5gm+aWrmr9ZH
Lw38y/p+KI+xqxH7/nYWW/oh7rsm6QRs2w7oqnU8Si9DOH/+Iet4YGVi5Lda6xfXBx4KBBhYKEFO
w1wAcXEceA4utADY/CfnR6OataUoQo3l0S82FuVI06Ev/hwMtpYYynWBwPhmiHOcGPSyYHOHJ7M/
P1WeuYpFC5IWUbNQmdtlFYvlU4db6eRVkPueRPbk2brUIQ5W9AG220h2e4dYObH8T1QUFuhEyR7f
sPGWvLii6WExsIsUD7yEWCa/J7D3gdVt/5jKFsleIL7K7+k9ElCVG4FfwgHpUQNyQfg9UIMT0EC9
yz7F1iU9pOvehSePL0/GMu6M5mIZqLSrH72He+i0IJ45/b2HoM03Q3F4Jh+b5Ws4mZwojhbYtWz/
JVF/ghOPkIChfiIoL3kjL7ZQMREb9xyTkowttjrkjiDUCiYefEewvVOTxqvlx4zqq4a10VPJW55G
eW5J+3fs34562EzQWFeSP5q6KGDgPTEOux20vEH3NoYQ2BJdg7v9fT19a70kVqjHwOskyURmcey5
Oo+nugnzpSeu84YaWA7fC6Xf4dpqFcP5LmfwYnvAfEBgF9VIpJlv/SApx45vYDShNM0y+SRPONAn
4HnOL+WCu5Lbggiqr0Wk7YPqmRzHT7NdtEKWAE5zpyCx10cEvMQMbTiDmYcu7bZWz9NaOxsZvF2k
vvY0IcCesXtTVBY2Kzesgxg1lS0CTjveY0XdYeNFyUMHiKq77QU1SQArW14mJYWCitdC2U/erZCR
3rzGChxagj7G+MyoijiMPMYButmSidEUoBp6OpzZ4GqUIM2aHTX0Tp2kLQVkRtLinnENp12vbni6
0vlLbwfSUW82xN/1JH5nZ3sGLBVNDdebGGV4/WGtSfR70GJqGghYuA3ZTU/olNTb7vVttI7egjKZ
NUjwzuq38cBxDBtgxTAxM5usYGZshX8gkwOiM6R5IM6r9mj/h9V4tUpuN0zCj5yrkMsrqqAmCqZJ
kqH+F0fz9iAkN13SOz1zy2le/el7UtPIJco1BzdylUFCKCC9OL9Wcx83sVNp2xfWVh2aRdR9Nz9q
Cit/QgGgx0Jp566PpL26qyaqbQgi8KsizHWSyRl2ayX+dOe4Bsxs6uXKQA/F/d7tP9HuMtXsusWy
D+rbUcjX0rumGf5V4Am1TjSvSOc1DZk3x/DehjdYoUG06hMmQxblIlDnB12PRfNnA6BR2Q2en2CG
FC4JP7Su9lif1HCWWcVzlrqkEqRZ8lfvX3Mf47qUoB83iI555HMxVA2UyXcul8d5kNrDKN0c8YBq
cMd5cw2ygjy2iAK5uOqs1UnXJyhfXRBNJkouk+LUrLoil6UYYlLG3h6sAjudcGP/AHJgaIuK3tu0
EZ+KBl7pxl2HQcTf9ixBq931QrCcbg4i0LSNRvaCYLRpr/6eT2fUEcDR4Tz16W9N19hnWAUvq/Np
eqgguc0GYfRdnLgcvPQKCvSgAXDMlF+yNDLdOlzo9kpH1+tzf6eTqRhk3lczY8z54Kbz54zRQFlc
+o2xVUc4bQVb7Q2/rlv5hL1RoHRPOsAohjdFNwPSWhswY5xySfqn9JZf+pvuXKHL1QrCy8+T9+w5
86eJ5+QPoeQHE0FqzX7NK/YyK0vo2R5W53QeEOURU16QBJMdQxnoaydZiGkPTUcBxUtYULw//uw5
1wGz61sk4FjW+OZeXL/zZ73JiISq300TWl13TzRDJdnCF2Yrv0/TosKcSlprikQA/RHgUdvfuXPA
pY3ZZVV3q0RtcjgxNOc3QSgI9J3nTin3mDRhnuURLwlYFEibz6AMEPGBj3tNy4nocj08W7QnZGwH
JNk6Xl3OLnJbEaYOVWjEwmNYe6R0wIb4RFhrtOSUqBFBJWBI15L/iC/tIpoPd+4U97MDZEnyLsfW
pfWQBZOH2gVdaOiekdnC9vPozRx5cYDnG2Enu89iyD1hG5D2e2WB1oLFINPDC3Pf8t9o/rkGshsI
3m/s4n637o1y7NWoKvrpVA33xnBpIwuYpD7x8n5QnVTHt7hKGpzEbjzRWwAJLRIqu06emDABZebT
bdPO0Pc4u774dfEKw0l6EnjicRisc7Z77kPm6Swwx2gnIKpsQLj/7kGcVX5Nk2SLcH34T8BFcsI2
BOallgAtcVsYxskSwrJGn+G24wKD8VovJ1BV+bhnNMvFKNkQk4IPkEza7kHFn3IZhRMQtBCiNsU9
EpGrJhhSqDe+SxnEvqaaAoAagJwbmKsFFf3Efr+7TL290niBGa43S4lW1vz4aZKYsynV/7Jp9sF9
18jRbddyI40gnxw4dvcumbbHkudu5VYWXx0oMMJI1RVSfwcgoTNT3un3xNtmMPKbPyejygPKQzjr
FIIhGVawmtFEsXjOYd4fsOS5xeXIWDAcyj/OgO+WlWHQVcFbNTeDUanTKVk2IQhVBP8BdUT7BBzO
Wqfh+PqLXQsoDVGThW9vAkubJHxRm3nK6pif8Y81BqQYvjPV1AIQ7h4MfBeyvpI4fcGRGStSVt3w
JpqDXX1wbtmhv4nix/XM1BgJ//ineaS4K3em6XJewcwJhmkD84hw7mfl/LN0fJ6NcSN7ytLw/BgK
1QWL+WwKGa3hlH5RcHDqXXh460C1yhYtR9Qf7+sk8vQQtv4f6SrMsmwfq5vIpt7Fq136+y+3qyj1
tGshAup1GS58JcCbA9JVAeBjIUq23iPuaJvdmAcOLsSlIUK3Ag1+a6h6E9n9pOw++NmzoQnaSaJM
nMQWaqgkty0ilMYvCFubZZN5coJmJ5PODd0+NAi49+dF7BVykzJB0nippOOxVEmM2XjHWsZC9T9r
zrDljaav7hbqBghkrJ1HDhM34ShNgRhQPlLx7KLmFn2uTNV10CnQAdHmJvUYCcmZXpukszBK7OQt
Db+1W2+ORsMk48N6clQ+08tCkc7J0pOYJFslHSKOVGS6EV+wkms1yJ2DAma9LZWF8q6DVPwNhJ9R
izEQyarPo8vco7XcAAK7ODW23CKslWmXjXjq47GJiucaZU8SYOQpSmIV/PYrFvszHR4ZULsBuixB
VhFAHmj6sCHrNDQG87oh2gvRbQ3MVrtoRvt8heLaBIAZCWa0bRyOelpREEXNBRTf/eaAH9bfgR6T
OtZwzQrhigw7YRwlVcIZjQ3EMZCEdkupyJwrK5RegA0VILII/LLuZqTA3+5fp0CZ3yyNlaDBq7mU
poCzyuq7rIfoHdqO7BR4RWbRp6uvB25Ie1uaiN4RGOwt/yVs6cvVLcLUNiQSx5iSNKyyMBwY51i6
82BkPTIZsYH53lDGv1hMPEgFpF83G1Wo16uSh96dLFjWpfUddGv+coIBRrLEZmrkdJuRnVuedyvX
oWf9doqQEDC7YrgSuKPjZaU5glN2KczA4cKccfgn2GeaSwlWIlMvc+rfwjIjDZ+zW91igt/TBXNW
eavLlkpHmoaGbdDIFtfSqPNwVA07Tb0gbwfzvdLRIVGPMvFJfjkG19G8GKm1EFltn32M1OJZX3II
Xqcp2wWZQNeAO11GghATcPz5ZwP8+rgRHnaobV2iKdqyAHYOdAjB1COsFOM929ADZMDrosGV1w17
5H3R9Gem4U1UXjnBYo67DhdeD0vMC4eNGQqZPXYbxkFLkUfbWb6RQ2qlvVA6mPiWYYkoCd7PkEo1
ARgHtRrqhl3xvKc8Ge9bgkJDmsyuxwfkwOdPjroeFIfSqXuyavLu9PCHUpXOEyOqJPe3TXPXzvET
tj/F4i3gpEunmR50qIGBuZ0TJjOPVWnpbytAhCgZ8qUFIA69UAQ15k4WxrwOJHE0C9nJXDmsFLWE
lRScIikV9mywBd+9JvKh7rUlYAfmybUiBu0BFLrP8INXW0SMSS7as45xSNgRVvZk7k+PVU21M7UG
L9cKi5pBCzDHc3rFxfpjJceJhisYWT9JIMH0CZwk6oNOLpbQh+6QUj0UFywejYS1cYdM5zVjEUN9
02fu9feOF5/1+LNGCXKlGrqCGBMwwcxx6oc+eLu0vbNuq8ENPAxR2gCqk4XtN/yg29umFR65LkHF
FKdE/XU2TNHybzNuejYLRr4O6fRNujL11xpiQS+KgTy66qxgdAGsPV5fxEumMt608a0OndsnYwBg
4NNeHJqpQtooc+kbzK+5yQQP81tvuGpI5VJwN+0y0tN6V0+FFgcL3js5hB3kStJayLF+blmeqtKD
e/Vj1C03tZPP54aymBHzboaPEtv1h2TWaiUE7wFGzjq13XWhLOM6PnRv8IAhnjaPrhxB5ZHHg9jc
pbZ4uJMgJcsUVDipYAKSEvKk/Q5OKADl851Dpk7PYkwy8EHJtwq6sqYMhq55Dx+7fLXEr4RVLTBh
RncRHQAKXLnWsBMHgm6dQsDhxdlYw57mtNYwBb94K/HqTGxeHxuYWOoBcvjSM/pkACqk2PrNYvEd
XfYDLVXPaiLuFmYtB3iBwoXlNk40K/f0DfpKf0x34yXSTn14bCL9AILv4Duhxgq2c+xmg8ZjqM/Z
KW5fBusCH0p8wDoDt07x07Bjm9vTp/K4HIRHUzZBkYH+bPh0OKAuzkQe3bYpKt6MIQXEf1nlams0
uc0QqIMBW2jahhSNHmNI0oL3GjQa+Yuva7eQ6fmdFNv+SBxmpKFIiIASLeGkwziooa6pQGsc6A07
9hln2bK74/fac6uZZuuMc95qpk+M0iLuanxRX9LVTeKcjJ2qx51w04Q/7ck7XrumQn2sB+vn//oa
BAMNynnKqh17+0YrKMcjnojOPhnIqFoTOZSVOYylx9xFyhb5aov1BcTFzuV3948S0Uk6JDvqxq0J
LHYtBfl00gIzRLiCsaIDoHOOiG0W1zwIbqErOZbvZIfbzLptYGXbsVMlhR+i1wbwRWcBWsHcIgzf
6zafvBVdHbRQ2J0bFe7v9xenTMbTA0+YRnxR4DFWhOcmM8LrGj+au4QXB43HV9fJ4Avx0h244CVy
k5pcdyCjLhbjGSqCOOU4wMsAKpv2lL3lfGzukPgWRH+iFDP2gnOfAca2p83ihSJ7P+SoX7tPzGNz
LeZP//dg+a8EDu+JqgQgF1HcX/6S7DxzMGWcoZUn5JI/XB/3UAbcjao0FE72piKiY7oDX2IcLt1J
p6U4GXgX5AaoqFGIU6TE/FiG1L3KqBAeNtiykfBdg54pyeMfUIExjm//9D69vCL4fGwz4oGk8iXz
8kIvrMDN1t314/YTHCNNeghvgfadvx7zz23vmEiaRbQn+g70kwms1UebFEpCous3KI6+aLNdvqFf
kPQoolpsOiqXKAofGx/JhZDXipO1L6GM6WhJyr5SQ8Xb9n9pfJfpGvD6polWAzzMtqfmfirbgrUi
z1Wj1qIFgI3FWfOcAWk6Mlw+U/D0FoMlxUBlJqahmBJLBzvxyJMJCBWjh5p8+7LQnEK/Gi7bvFc4
zLLwu5fN2gpKyJgHOzndB/j5D2avv1DZwlsRXWBQpal08/WUYZEiLBA5oORjZRIZNweiRk9X+SvB
V415ImsJnGFUSDmzx4HW14IGJrcwxCF8rW+zwB+oFDifZ0xQBybZPfLtyThvovVz+7HUHqXVGGKq
SSqS9yXmQUKqYCF8tin9UTBAQvDa8iVDyoDCfS1OZE/O8zHmqrd0CRGF6IneVa1jiExhP11Qskv8
Sgcb24f+SfIOStmren/WFH9TBAyXmKp29bjTpQkm/U3FdzJokZ1nitoGyjzkUZSCGv/qnFwmX5jV
UONWsMuDfR9MRyr5aMBhLQITiLpkgwRaw8Q8AkmahX5QbwkSIgU+IWhfn2XwBVh9h/3K2FKMpZ4f
mT1AXxgpTRBizY48qRmCX3MiLi6+pfjOVz6bljOgNIrNRAnePvv4CWRYTbCAxv/CaM+6FTEWPTOU
tFkmbMAbiLLhOT+29f53wiZ/537jdWVAZr0fYVUhu8LN/qI9v3noy0/j7k7Bm/kQjdSSZS8N1C4h
sx2uccMgQZQ6fwVhycHBWmASeSfl9bMFDYAY4rd2+xzMr6Ty76bp+DO+MqKPrbJiS78XiKAj8IHN
fKMT6sRdnpzWAY1r8BE/4I/FcmgWtfNHPX3IbbbI6J2rvmB5IL1dHB7Y21jXoDPaAZyqPuhpX7g2
v/vcngCJQlOhXEZ2h0uO7jrW3XDrWJhTJc2m9JBMjs2eYvPEoMslitMvQyleLPPbgPnBaBpbNIcV
KEjcc6wnaRJjPQh8QimRYQj+1j/qy8EtbmzO7M1KT7nbtuTSS1VD6+d6KOTN6jBcG5hNOdekexjy
soXE1cDOM2pMXLIc4dUG8Kplw3SMmj3w71ra1KeVJH7CIACmfMoLHT6GbPE9A5KSEDBhhWzmkNFK
7Ydl1JUjJVggQemiqHMJL68ymED0+LIon6IyjOshek3GMEpkzG4Ls1GCEvVIDSxG1iuiunTNu0/K
KTr9yUpZjZcN61IZ68mHbXnaKS71m12ZmGWiItkuDu1TOnsDKryyvjmcO+Kz4bBrS2ZJJzHCFvW5
5cuJlKGJ62GPIRfrRWseLnEJTopgh9QwNSmKLm9njNQpX7WAK73DqqVciMi3oa0jN+k8VY+qJ2ZP
8wtkfptcCPUryOPcggPWjdDK0spGmNLdhmpdAU8jd+j9bE4XmzPHEzqW1QavHiwGwVdgpjt3NOYc
9s3OeskWGUqKq91R6dwqOUa3L76d12qth2oJRGqR6Hh2JkwOYZKVUuGqongSOv7Q8sEqUcjlEau2
kR9dLr5OHCgluK/sBvk5HBzir3F6U+4qCBMhEv5LcjIKpbIa82/P123JfJhSOkIbg9CkO2S6cpXu
YhQx+cHTBdxqzzxG/3OvQ13H+7rj2W9gcZOdGACYpzETdSAgcKLsHzjyk9HxCc4Dbz/Lx0FMuXea
YERdDt1bH9uhVwHZ/IGVjoT0awDhJUMhWTAQavx/xSNdxqK6Y3i1RPXrJj4+thIM+FMPSCdiBz5W
Nad9QX1ca3o6osOWzdc7hiCFO3QB7R2iwcOhR27mCpRffRk4+z4K+1cZkycINFDt68cb5pEUlGU5
EY8kOtzNO6HwqnH38ic6gqjP/h02YlqmdB8WTr3oFF94RaVQXOZmhU6J25ufolFa3+yPOa88LRW0
xoji6eq+0dS4LhuoOvTWPMwkO6C7KDkLYrUKXTUGZn5N6ETqs6FtL9xQJYNs1/bAcqttDHuRhST9
Ea1OlNWOOCJIT0Sh7HgnijgfxLmnxG75T4bpqt80farkuYWIUfyL8IOQXHNxRIAxfAWEAZzNwvLl
x/k06sEgSdbovevtCl/rsPl+X4iH5gQWk2sgY3q1qydVi/RuC1I6h75jYtbdpjJyZelmguWmoD85
7KSBLEdXORcFxZ5HcSSniD/td4jiGxmWZXPagFGEcIByhAcBIfszUATZBPKbfyxRd9aJ41NAyxTe
+dCZNzih7LEhacujSFHfSUS7znVQi/QobkmCzvJu34RfI/P5XuA79F9ApD1yVZKOrW6QhwrhmCue
YRhxyK45HbebfFWOy70wscnj+PnSi5IbZiwSvbLtujjpQ8lEQojVE0dJ7eFN/hQXx//CRLzatFgY
KMlUHXkctLJ8l2X5qRiBIWD0dtJhObCaOdLCNOIYTaoETBWSkJWUgAmGpjhcdeP+d4C+/j0ZxJ8b
mGfh5tGctsRZEH0yZCFFgRpLiRQV32QEB41jTwvZ8l5+8Voy1Gw4Lr2w1HzHwX0wQbxSKrzR2ada
BP6Nwy0eBX2jFpL2KJsu/YqD29OtX+TTXwEHLhJx+dUsajIyeSyjpXcrjI2hBRR2jXYe9m8vBXqx
bY/EC+1SZLWfigs8yBWvFml4W+QlIKc4NhVDmFiBC3vWlqLmSw360oiDpGWpz6Y5iCc2VeUP5Vwf
7eWQALg6YpgHeyxbVQ8sTwlkCFLM0Tz2X4U44K+OeZnOYSXDDdHIdHQ1a8L24B0fihaZcNdTVk85
fBTlqOsuEFRK7eMWE9CvlmrKHVFDZX41/qg2VAGQCKLcZAsVGWfiHUP/eWociiMzZNw5UkqKYEcA
tFzHEsIaTKVAhKeDZNfclQ3BBpNZXutP9GW19iOhLQpFCce36G7nvpkrfYE5foV13kiE6FzpinrH
tBrj/4KZEgMsTzCcnxXoG0xEFHB2ZvrbRfrGdUUrvbP9vjxU2ymh1iROxSPkGz1PQFYyDkEs8xAV
4MWy6Brt+PuacN3CUmBUNSQ4uWA8EOHnjiFyAo3xK73u18QgMPhPTFV7XQvEcAWyYyXVcGk9P01r
JyX6khdTN41l83PotZPyLf1F7N03jwTwKiA9Y7OymXxPs9mMbRrA7o9451xzVEc4AH19lfS8heAh
zEz/CktnRa4djWXf8aKXb6sWtmZ4aoe0A83C68OdCIfJx2pmkTkQOvSsR6G7DNnDgPfN+hb4ngCJ
x0CWt84cM29lBFFELP5AXeDpYnmj36NHVT/rNQIcMVGcSBGfqiWHAgmMB8po0H5yScRMonhpYQIV
IOUCeiUrFg32ANDDN45IesKylaS19aJi6++1Q6lHCxoTvj9vxuMMrv3Sx4x4v7ZAVllOonT41k9x
8VNzdj1EtAv8S/Uj9tYvvJf5xrsR8aFguuNs9jYe1INCrCE4tgLC1OkizSqkWEyfX+QyhlCfRwzo
4R6uHFFbkI8CYZEB2DlgqbW4vjg+ZfiGzHeUNuN+AW/FF0iOKvE9Es42Dwdar5cvRgIvcjyhXuBv
vP16zXkhXIkFYHg28jnpXhlZJnsIz94FIdTq6DqmGUHCuSUlJpe4zCWjUFfwgbRFXbAcx44ybefB
1kcELfauer3O2WJrp3Z+sMJY86ft+7seB/WMQ28dROEM9srxwu5yRKZDqUIyORQA+RtV2+xeKS+n
Z6a7t79dxIDx4LjSrBYVjWw+D//Z4/HTlm5KXBrVfZpgI9tcoVYznpQ38SlNtc7WcqGoEgTaxEZ2
E5AXX9HQZ/t34NPWB5bZQey3amg12m4GCDLmgiCT2rt0craAb7BmYKuIvO3AHd6pxLnqUr881gPq
eSSYjwtjULik5biDLtmJxzgDaYzoP1JtvC0lf19h4UdSsXpQaxsPRg0QHb+BrkkkMwBdR+9eNEtV
DKfNKs4Rmc6EEHsOL2k5Qk8jGthSi2q6s/S+RkXQaFjBhsyrDaItrVdy4SkH7JoYD6aUdw9KIeAb
oqEPWUrKjPd11M6nHdyZIcdz0mr2UVqumiLLHp6LG7GDv3kaNtTVzr2en90/lFSIyTfS3buWUKsu
AoHiCF0F3a1Yy6MfRiiNC1pskY/7hA0oTzRFB7vHqjNKqnWACDdjrHzGepXRFYb0pcworIN4wAqQ
BqXl4bn+qPBfgGM1SH3X3P9wygb3vxS50O/1gphsAzTwxALPac2TbV9MsgxLtmXIxHn/LFoTes98
I/pcCj5YestVdidlIfJziU8aZPpArmMNPiiKIRtBp5IEooUqD8RzqldSdQzcUlDzye9ZVZW4PKym
91q2DMofL2FG93dnT9FV7Zq8e23B9GhuR/cpe8r4T7oLDQCoUkSgDJfPAPXE/jjjLclsBgKwCrO/
zvFHKtXgi3+ULX2Z/aRa+/3nRVK/jYO4XdvucTXXLCgDjf9mMpUg+6f0lSYoUTeVsBI/0ZRi0kQN
R9RLudbSsqnTZc6LAviTr0NDwrVFTzPMjhxZ0ZvJPw2syS4zE/TeoSkNC2777MPPqAbo427TbRSN
WdOZXlWv14PR/zLUri9w94BXXMLqBf5MM354ihSoFrerCKqg8cZKz9nF0YcKn0h7DZr15lwmm0Es
khKBy+PWo6YgBddRan4N9ujIwtkm3svbDnJXrCVufYv/tm9SmRCMNjyB64Z2+kJpAYNFgL5y0B5A
m08qnhwQEnvBLZq+RNHAACwHX1iaUiIG9J+lKST3j6wD33nmjSSf2W4jnMsJEOfuaU6uvOgSPA2I
X+UCkGWWRTCIZsTRGJf20USNLeWkPA+mBXzb3Tg4Badm22bq9QLxfh81E9Yn7FNF+sT/ppAGNzQr
k09qYpSKaPx+5TlELU5e2XZ8K7YGJexTtXyNck6QcffT+4mbc9AidD5bWL0a2wy7zYRCvHPJriGq
v+gjXKwS2ke8L2KjEuJ29eciJE0RYs/PPS93Kcykd6a5m3XOkfC6B5pmB6Aqp0FRLT35PIE59lpd
NEw6Bw5qa4J43euBAlv2CimOTWzAH2n2d7v25ObmHR0hMNvzrQJuUq9lR8KFsojQcNh9rLPS4NM5
aZteUXwaWIGwtdlcpeFsrs22UL4SsTgv35NyE4LyQ4cjgKmkGoevTrSPPfw6eC2yJOtZYZcMBTng
S0NpmNlovPCwZ6Zsn2WaCKdcsA+iYPN9A3yvAglG4e1KyeT8viGXnKRLgRdBSEObFbfJ1tbD230t
8dE+6VrEKVwmHx2om0nqzc9zD8Ibt0htGMfG/k/+veTQmy6kzYB15y3P17Z6kO24zpNopZYEACAt
llOc+zSj5kPdoS6aAKK5PjuouMzr1UmcYLlftXnir192R//cscnVQM/nkcXE771UyIwWqmwaU7bY
tkRx3k+qzJwTo26U7y1TCza3wNuixhr2IDJK8SkBx+T7IP6Sgsx1m2mVUlfgkSD0l3K+NkabdpVD
crc49lvtPFJZkgO4q1YFH+yxP8pOQYfhQKVyzXvwaeU5d0xsoj7UbEM70zUQ8OiJS6D7LBhn+oaN
4TdbHQaHTFmrAcyi65nENTpJVQGWKtY7gHLWmiW+DN28qRWQT+jL82TrrNmCX4CNcUKI+AdQbEH+
d0bdTi/XhzsIBTvD8GS9dFPONS/birpdE2eNoQEd38BdJiXK3GeGAu9XIWkJ63frOZ8BDX+seXKG
3p+gSU1vDQsqPHG0EdaJ2973pBl+aM1pbjJvXPdalOXzrMq5Uu9GwyMRo+fytJeprJcSV5q5cDso
fnPC5TZYn63HtgbhZIXI/CQWVcBsiqnAvuli0POG5+xGr4AMZ6EaPXo77E/tvh0EdxEghDwHN/YU
tVOlVnlG3uJS/KmjSoVwYP80S32Uv321lZDMA+nSWF7S9R5x9F41pOpE/lkrpOrn5bmaqdhNlyjg
M6oSAKYVQKgfvCQcDusQFM1J8dbRPHtTEdRRdlxjoUt05H0vRE9GVw0Bvhu0dLgHadabCSS9fD6L
7D6cBHyjVWn5tNAl5/WVKb7pYdOM/ejl6Jzjep27CtqEkNzCZ61ekVVt4f9DFFFnn5q201OnMeaT
HWB9EoDFAcMZCmYwVHmyak2FOADN4kTFxM46BzwyNhxm+IVk/keU8tJmaUCsvY8lJFVjOoRTEsde
TUa26APx071pEqUcGrjxOl7R3xZg4+gsXcQ1Lty/RiaD/txEQYtU7q73Jz6NpGX/qLA/X7Zv/cL7
+YVkyRRmDkIhM4mzno23Xg0K0vS+7ZHWPJBTQMK4af2Ck2esmdhJ7tW2gSZzFsVoRFYpQMaeGL95
ewGeHl+5A7YejTA+2OKAl3v/x8Gflskac3CYmOrCLBdQX/x3mYaAtgpWWnfWFBkwED+dRgw8DdY4
RIBKhMGFQNJ3ygSukwBtR+es5u4sIur51zv8B0CvJb5NiLFPaL8TchbtsOiVTnWtKms2ZQ+FsFh/
AuNdnmotdPb5f6OhcGd00dn+RJWIkkl4vJI57/c7AODy6HHWtRDKztdV86ZwKHI4rednKmrWZsCv
BxhnO8iu+CIUxry6u5obRrVCBXs1ILk/WvdjUEF1N1YE3HY+ilTXCsRkTovfSOxZjAF4yna8J1Pf
YCAQ2yF7cfMBtaobVFRmNl5MrS/UJvtlLHi60W3zYuZYiR/VuL4CVOBS6O8h35WBqS728E2dRd1S
rWk2hoXq7KqrWBEioEXebiqAg5NENpOD6jGfO9gfl5+UfL+kbl3t6VsAO49xGZb+r2JRE92NQyiu
oZR0VY0OUj40N15Wka1tRz//gnNcGEx5lR0dwCR9QWvNTFpIeUtvG1qxvAj2fXV+XsFrihECxBFZ
AX+TAJf2gm98gZk8Gtso/LcGvKoaRuA+wXAJrJcGNQ7l5xgWDZjCEnk7atzbMC6C8xuVtizE/pnd
bElPTLpi5onRq5Om3nJISNB6RMYx6FoA2r/MavPqEFl3x4tczEXrDLJEQogiJ1ppq82pxJESvTZg
JelScLz4B/v4UPszn+GyxI2iajOXEAueHgIkErjr03A9QWiYA4u/O7pNpke4GdPWK4XEZJzvmOJR
m1KtRXqdsWY3JuFMCrAWHB+62b6w9x43vvDGISzT7K6eMJxwtL49BbQi5zAHF8imovDoMnISusBt
TtTvX4LEzquSxa2Oj7PUfTkhTMRXVa6L7uecVWTmRPCjZTrjIqbZScol5a2dA5XaDxK6Tm8QP5vC
/S1Z20EgRwoi/xS45jzRRGV4gbW6yWlJYnMBHAwKlH2JMHkGXbeOjxaAbv1P1gesTSD1Gh4jYP8k
Fs4/V/FBSrdFqNCn+D/BK0CuUUkumq4Wrr1dufjF3efFA4INn5Qqm+5WoWUo6ghKylBYrmWMaJK8
oM9KfTIQbvbAKhIvFAvESLLwDP8qE9fl2pnzrUNiUGFhaZk1+eGQqGygOtv6x/oJOvgyGz14GCbL
taQhCexGEzks6BySw1Uunl6c0ao9e8mqe8n2QWOI3BunvD9yRxv+MLv6Q5Sc5nyk6vwq7c9k4+jx
2lh3x7ygBK9utMPXjhC/5tUZx67+YrQjr9RUikzC6S9m8Sj6CS34xi4ZtA+GDL6WOdRSrSDZJbj5
mh3kz543xQt0UczJfGUY11No4eNj8l0ro3wMWHPe6Q7ELeGk0ECrnk9tMHk5OyVUEHzeCcu32gXP
/pjnv8QIerpVPUquzd9DEDxzJ1f+fOwAm9HTDKw02+A+KanHaEFfwiDUEZ/LW+8io8xgAy/kU5Kj
L4S2ojaT9HWUdzy45XA7fhjJI0Sau2m6pDJnW/lD1u1eGqUGZL7f2iF1oDG7/lETnpxgj4dyQPGU
mQVk2eh/h5leIPzieUdDWD3/vzOySBI9vLT84F45NDQ1iW9atPkoc9mJN4oVpcgXSwVy+B0TKY8A
jK0nERAAw1P7blVLxq0nI2F+g0rKJ68VQe7i0iCCpyzPvsHMQ66/nmmzr5B0heACs32699Z22FIa
B4f9iek5lS7jRLw+Ha1Aod91LKvzcvAvsbVFAzFz2KFhKiJg09yvqlyA+4fVycp79aYeXrojJG/T
e/tIpcH5CKofvO++v2JYXvfKmOolR5WY2b0IFaXFwXkGhAZn18szvJd6Q97wbt2OXK95vYaqo7HK
HkiW4xfpqGgZK7rWol0JeryY5Gs7r2OxZdL+2WUIAAubA9saF7EyNYLMwk2mFsJKsljdo6wrxNJG
+bA51BolaVsLYLo2Jac3Ef3HQTrkQdkulsHw6EOIezJMGJHJYHzK3SgNSJ23p+rrqHjTpAL+HS9c
j/09UcPNPp6yUguuZ0B7ytACVi4ZS5P1NOYBzg8hV1cF9HF/qp3vPyaOAcpvfglnpoO9hOoGSE+f
3bmwbljUaUgthxgK/UTkD+L/dl8wwbvN2H/iOs1X4qQKp9axRA0mjjWRZpYfTyyqhS/SAI2fhM+M
ZVaBM4aF3+lzTgvNP8eGxUeq42otliMS0EX91ewpiToZt5pJZ5CISYNBrYvltp/hp3vvST0LykNH
56ytiZvLlnwC0dJPo1BmGZVGV/FLmIRq7eGtiYM23W2e2E3b/kQwIUyHB4rSJcaPxfBrYBAAiRT7
lFXRVWgRftXD3cAj138nyU3bvb5QsNMYdgEGIMGt8bKTr8HXHcn7iWTYKpZkut5nygQ4wv6kxBOl
oOaxp8Mio4wcMPBxpYGvioeQRef+cN39aAjDa+d/a7gL8c/4oKgakaXM1S1FF0aT/y8Cy86rwITV
315iCsLcO87sMYQ3ktPkUrdbIUF6IDXM5JMaLMM0O4H5wYXBFXgUprCagOx0zCCtXVKLY1CZ9a85
QJx4tuYSaZgGEXwdmaEMtG7Q90fyNVLKYddo1n5CpndHohaBubDf7HetSYDAq4H9/nKrxpmCBWmQ
uAaGBxCzIBPAud4eumGCkYjJHT9wx1ei3FfAs5w4HtT2z/ZwkYXfRZ1XTmbaVULq+61R/KpYANMq
GtViySeTkV5VBGUza1d/mhtDupB5xRkHwCZ/vg9tjCn6oh/uPI5gFD1fk91vlRCbGCANyPYmscYZ
xCcKa62rCXhZjpUc3pk84oqRlEFnIYhfsF32FQKsEWFkhY0iUtbCtWaBZxeqSDDieVYUZ5Uj2Bzk
nFb4AfrwtvzinlE37rhFgviJEeVBvKdIO9Bns50juOnVvROQ67c6zNjQVrWmWI077DWlZS9zz6dX
XSGxgvxdkNHMojEdva+XnwcvFFVKBJFXBTyS7uEo5RUbSA40tDCPpbxv6QUfSlbhgzpk4BwacmnR
PMflJ0EvrUkZEjP3p8lsR2Q3l5S6rE0bncbSWfgxVTgAdFixk9fnAPGzmAW5aBTXD/UNcn8q7RgY
YP11/Oja7auoi/nOAWygjmskDD6a6hcOLTHftI6S2oDYm+dRHbG0KUxsrHCBzKr3QvfcnkXVRwVF
00Tjnd6wuftRCcWbVm96ho4j6YCxe2c5J6U+c+LX0xltfac5Wxkd2rKQTE5g+W2Pz0knyOMA286U
mViw03VcCeMWp45LYM0G9Pvp5XmR22veI7UNFz0PFh1tzmXLxBlaEVu7/ucoeoZUkBXrkb2tJmTK
oIBa6kIpbrCy9GgjefVpgkRCVMtfZJ4OqVea1wVcONQ90KdNLahKqPIHFYZpjExJcgTgA9cbSAtM
pimqQ9Fy4b6xMZD0TcIW0vISWrAhB8DLf2Re+C9xjVBeaHQAF7tomPTMtb1YgEvFdxzgJJcnsCbo
4YukGYk9/RbiabpYN5HYAnbaKE2GHmJDVUNtuN+q3S2cns0Gnigw/Q3Mi+n/TIMsc0aTfiAf8SDb
zyThrUowsqUz7KOQDpNjngYmr1Joscx6E3CJ1ePTMQLZGaKDPCkMMjmMbZ1KdfnpgHuCTgoTk+Me
Q6CQTh1Vx3/m8fo96iIn40WJsEzdIPxs9V4CMMv/uiPoV3VQmsyLoEzYBii4RMnP/u/RBbmsHCk7
9ApCPMQ49tp87h4wskCWSl9rQjIaCaB3OA1j0Od+sNa9TbMAhLza5rFVysoj8d6NbAVc97zI0POs
+a41WFJtjFwFy5yV3KBna/1jZtB1GGpv6aNjD0MPf0UEkD9aRTcL0idyj/zvs8Ls1whlFBOvW3xV
yVRHiz8Bw9sjkJfeDgWggjGakb5W3E0ZAw+180f+dnELhjXm+aNkn+T6RE6OUx9kk9wfyHIEhn+M
yShE4a378lY12UkcZA5uvwvz+6krnzoW0URWPeudHPZNVYXLAh8MKooj/+5noGwS+kJVCNTtNnkV
chqK6QmZKGwumo7M69dltsNeMSflwvEK6RYlxcCwFqxM2CFfle9nCiyfrOb0U/qxwNGqUrTNFyuv
b2JmwCWowfHL8Z/MkdBuipZU6HwYsG1r1+UxSnrnM3GrYK7rebqoqmWrz9bLzWaTwzIqEDP+qDXT
FtLQBWOyBuEHU0Daw9bAZyAsc794nJ8AgEizGqRd73vWe+KYgQrd3h96Hw2VplO4t0NsgIon0+vc
+I+eKq/fKwPDV11H5kTjeAmg5mZtYntCp2RwSxYdPSxEH7vTgV4JsNVzKzFIOHlGK/aG3HPg9DJf
OXJHijY8aPulAtou/D41X+8k/TXopkYzXbYDTbIpV/ViWGKVBsXxVgdm85klbRodnFSlgtn+BuVH
cOtOteq274lhisdgRv2i/URs+QgPsRmNb7P1hxvnn1/01hbyZIVTdLbIW86ccOwChcxGawNWxnRV
QQN1GtvuqgdtuYJgpUhRGwR0X43AKRd7wTtL/UCYC86JHeDKnO934hxwje3jfLkgjnGeJMn/1LBu
dL7j6WhOuPBL5G+KhsHinWA2Cz0LYH2/EREe74uuYM1rWvI/XPDwBwEDD8edTwWM7DEc6KXb0oSD
6UmOZb7i3tklZ258nkoLXAqGhCucgzCzC0qp7X9LRG8PFUAH3FgVVkQM0Vm64f93w2AcVfSiAyad
FLvruN51aDYK7kxzFWFurgg18JeJxcn/mnYsCW9MzPkhMpTDNGgiiPk2lMlw8aVfyuM418BdJySo
28lLG0qeJy8OMbzMyZ09ojjTxGw7/uE50zF9IZl7++OTsKuTE3qvaxSbBRdgp2jfo+xEbRtDi5e6
2/W0wxcCZW8gl0zBfDgfy7swOeTGBetdWW+p2H0Gl0J5GPgr/VVQXzHC1fwRcTe0uk0C8zq+3zh5
Ss55FqCE0YQuUAjkchzdsWDFz44zqHnvZ94IFZpXcCYpZ8Yf7PGeAL9Bz59OEuQ81iBSSMIhsmjp
4qRR5Ukfqm6A97jUiEEFf6KGh5qRTdFTg4KznZAx421hYI1OmPwVjCnPJHP/i2GNnGYnBezHptVK
bHRBDDQ6ebTH9EpsnwqHip4u9b7zhk+gMhU3j66Mk8sskSTCMaLty1ONSLocIU99HzTcFFSAPUUw
z3SdP48jU2w7l+l8VYzG5ADfgLHvkc6hAI2+0V84Fwjm7uHLZGevhn6AitVvbHWMgfhNPuOj04W0
bXc3KBxH8JZFViiBxLWjAyU0o4rwJOUJc0OEY136bfqgMCxPIJzxSFE7SaHsvtOZOV5CHVsKXc0A
sLb1UarFDH0/0ez0C8POKhE5XMZL/zx3HgxxBQkXRP/4tdH0fJfGR6LiquFevMW3ZtSzlfzPVHr+
RmA5VEDEkufNfMMnFQw2PLsaDpqKa82QHlSEPpNHK8HUk2lS0aw4oqBVbhvNHONHzcNxHvIW2pNO
wSD8xiCKK92ketyivozdCT9QJstEMEcR3O2WtvFaCS97xXZZIhhH3rzPryFEth+1YtXVZf6Q2k3g
SRXae+9eOiuqUTW3+ragzfQuKtNfB9+gdzm+tQTSLEIvUxLxqVrt/d/9srbZxbf6BIcpzJdAN/Lz
mnOFo6qIJ4ZqhKyZsfNO/1/Z9QjXpd7/pAOG3OAECsS0wPgAZYzfjl4nK2AbQRXe5lK6WM8IN4zq
6KmEOXKtWqpS6SdWV0iQb/Z7IEs5EelmnNtgjr1HC7cbi74g9lmw4QeN2/zzWFx97uBdbkYoiZv4
vY4UIU4yDHGBb9qFcECSb1yyws5ie/LpWQ7jmTyc4ESpOiDPf4ypOTAxsIhWAicddn0g77xENNwY
Q0IkINFMVvVv+ZleuJwQHynnYcrKNlKL99+zeI0NaeJIINQ1vg6GBfH8j5MSMWi3P12Q86KYCwiR
Rmd1n3xx9ZkTCpgANiigFcL+mvNjzYKwjbu8w8tSi+RDNAFAHDN02i5ChDlZgUv87OtMqYwPt21y
FvDWoKrb2lDI7LLENVMksn/BVlFH3KC/+1XNIzU4MQNGruk7PT+uxAJ+iEbx9i+WbevRMWzZiCLH
WTXvEN865S4qJ3p5szkbnEUgJkWfg5lA0TLeZu33zwHdXsJxIfkiQhGcqA2I7HD8OiyXSRqnjDVW
USVtEhnTEoRD+ghGHWmSJbspe0J9jlhXISlPp8c65MEfkveQCC7yxLlqmZbYG4JeBI6bnMljv0pv
eFinB2fYrss22cZRbfejcUa3gjuN9oh5b2Z6OSRRiIbM0qe1lyghJ0wKdnxVNI5S1aMLlMZ8Vk/Y
j8UWmM7RiY4WwgJntfk7g5X7Uh/71TaEjTlYjp451bNaQI5/MtMyiq5oceAjXEXPJwGI/AKdzjeV
TiAu3k4Gq3LRhoTr7lH+0z4xXr2drHYjzy5ImlZcRDnEXXmNWzl+LdIlYM7T30/AUgTU2YN/gfoN
HTOxHhNCO/AnyizoGjltwOa5AFtwVHwnKsAOYNP23PZ6choBdAI/CZj/QFyHgz21McT5jF60ZQfi
8flaUef5zIbnCXPFttaiJW0eYHccL34+/l6YR3yZzp+5pmymxQiNr1cP1XIW28z0QoIYqQD33oQx
+HASOx8RwUivZc/GH8xyda9vlKy1dfz8QT8LfrmTQy41b9MPkhZFBMooNO7CdlixYX/Q1V036Blw
YgC9mcWkZeHvz5ePgs7mh7Upi33wsjH12dQ8Xsirup0xHBbsS1/w81tiYsxHQXvkxylUcsoqjP+C
22H/ctbPcqpUqu/WxNzdY6++47AW4E2X29SfXyQYJY4wCzzQ51mOsVivqVGKJb2Ip/Bx9ua+EL3D
PJQC2TIGdpy5qwf5Y49fS9+sW+YlghJayFvfgTTD8GO/AWUzid/YDcNi4qrXKa2u/nxFdtjHIBio
3jHtwnKeLMyRhy/kpvgZM1h9LrSX74mHloIjqQAeEiecnn2UiijaI0ugreQwITg/tq+CWzbmWHcX
BEVaPWsuAfQxPMiMVrSUjQUB9PwHO+VR2+wFGrzGwXMaYK5Bmgai8XQUCtawryklS/fko9y8CxLH
SJ2GSp7vzyZGzW56g64btwPMtT74e4jOLP7B5fLywQ0nJzCwyAiqqU6++PhkO0QmzyE4agPQvh5O
vwc07tR7hdczkr9PEmOUtRKJWC/ilSgIYj6R1LLUOOMZzpFC0Qvv/2tDisbDvT3OrVM9iNGLUt02
oX2MHVR5Yk9dxQMiscQ43EIS3QzIjXA4XBGezTGC583IubdoXwx/sLysTzgTyhiaSbZ8KUcsBErb
p/HncS3q3xdkCX0qoBmRxUcPK2KHq35XdJI6NscQerVG/im7IAmcJS+nzraLWrZEs4rDtlvvSuD/
6VCQ5LUPBaFrPcJicbiyyDITSeC5pkkAbOkmdQsbZ4hqcEqWIKDPeSIY6Yikb2Ps/i89RR14mukg
udceDnUp63kJSViC1eXPpEgbcEwNTD4RizDSTN0hhyAFXJ+/MGYeWQin1wR0Mfzz+mTH1lmQflWd
PNasfZiugDqBKHp0RPRhX6o8MIv8RiO9DfXhipRbTrP53W1GeCZ+D4xRkbG5Ujvq0I19lZlMorR9
BaXP/+3h0txGDsxk1IA/qL8W7VYS2DBHJY3FM8dm5B57zcVg3mOiIjKKnhUyeXCG/AypTE/m+f0g
/RnIVRmjp4FNTGVOi3vG1zTwjKLAZq5eRj87+knZFfptTWRrUJUGgjgEDBNbd0RCdn4GhqdzwOfR
awhpV6Cte9p06oXHjKQ+y0P4x5hkUG0LSMkwhkZbGqD86XN464CskL5/6LHFuXWISjlX5MPYwx2M
5m1ViHlFMKD88JQH58cR1ty4g94Vhl7L6MM51Hy3Hzf7tBfZbZ9lpLNoi+KJvI4hODkTVCP0Tf6g
98ce03YnM7qd5A+Q5O3lkqVJpRe23Lmm0ewz0dHnKloyEeX/h+o8YpBxV3oDHqNwOf0erd09fNCp
ZW5rsww/Z8Zz8OzZS2D6Tsy2chesWMlru1t5xvnm6/UryW2UbKJkGkx6W2HDmafYMms92PrUAbea
clg/2gllA0Ds92jgWPZuhqoCoTk55DSP/fypz8x5IDFznl2y1R0/WCes0Atm0jWpW8kLFDUjlJ39
PhrjI5/Htg2Xl0YL620tcHfNEF1xsbRDa9bPare6oMxN/KVO6yPGpB18Nybk71SmvfPU1O9NIHhD
hbbizyWvz09+/lB5Jx1eBZjDcj05CSlWvCHRNIEYguSLyUog8CbIqHLpLngVDkcJKpPHXhQKa4Zo
dYsN7TpUVLMwASBcpChRjOkxFpz9ZC9+b/xzwZGM3POS/eYf4trWBs29gxC8ZzbzIUZkvk5lGYdJ
zjuv3qPZGJwheQE9gV8f52mk5hhU9Yog9QOxW4e0Q2tuqTmPIsjzl6aaaF6KBtl6rCG8DwCfnjSR
KEsUwGxGeIjPTlhGsI4p19KcTRyv2pMu/ktB1GG3n6jfQdhUcDbcyUgq+zjtlhPs9pfm+kNWu2MT
AbVFSeO2Kn4JGxwz700cW0CR8PzLT+JQBAwpMSAiXaZ6FDBFBqqLgYCiY5tcoaUlvpv8My/kHv9J
PN362HplZwJi9Yeojyb2TZ2QB8u10fuJ1YSfH3GZ8WzSgtEGc/3hSxzqNsrVPNRzPIQVDCiEvVEb
tsOwfDeJDGSnWhz8SE5sMkaGNVbPB1z7aAfuysh4W2soGvgPRp6wDYHTez7bluH0cQnvAzjoKP1O
fEGOwOegsTYc3leOaoV+1Zn50v3YWRguANUfjgyyds2F8PipKiYyjoOBL2p9aZVHR6u30uwgdxCt
G7tDpbh1YI/KIPQv83AXAihAHV1eQ7afkLf9rxR9opO1HKAc7IoGXfRprC61letyjLkPIaqwLUWz
HapRr4w6ZWLGZxvqxfPdP1achnZP6IOI9BW+zBGjHzll6cz5m3Ge8ItUfthioryAtwIIMeKOajlj
8gyokpJTqY4R5NPxzxWvGmu9A9L+d0L0ENUUojfdnhL/Z6M9rwNCncMel7PDZ6pbxCczMU+KKGsC
z4/kuOvN46vngiyVjF3eXYa6fTZvqm3lgnOZEnbMY8hBpoo/AP034/MBVH+4n/TwG+0IpHvoItBI
sGCMmmG4qvlk8eWlYhCFunUOx+JIdRW0lamTKAga7IF7tYfFyNB9hicMSuX1B+xrtW2c6jk0dTPj
DP8I7WHLUpaBm5CQtPEK1X4BC8Sj3TkzPzAtzjv42XFg9jGxHeYg5AuDAgsmTW6UUaayys+cIrx+
btDgRl33Xdi5WH/1fiWZNB3ydebS026n8KM/rmRwmA+qlMaGZ8gSN0FkiZXqIuscdThh/OVmB1TZ
AF6q3yy8pYT0XQlM1lBJ677mdkeDv352KfM3a0U/2b+/rhZqlJZxjlHyZ0koJASamE0yaVVbmhzY
dPBzOp7iRznjO9yT9OJiVjoPrPi0X/qhTaz5DZgl0g9tEji6ifHeH9qdlR7DlIar42liupx90Q0x
FcXrl8DAaoENRkhg+V82B8WAp/9mGvyWG1Hgi0HbRCe2Xy6UGil8O1cpluSWlWMbtzlVwKJ2VE87
GGTQ1x2DOuP3SXkt8/jq4cDdUPXkucMybDX/1AaiQ3wvvntyDadfkscnxD/qwWSVVHeBXTCD4Zli
KTWOcKlkQwXvO1ETAX4Lp1QXlwb8xArK1d12CNblFMiWn21psLG0TELpwDI1/MTtdJFNYwdTWup+
NkdSW8bqDL3TgTnGg0P4/VPh1losEJCXKh37/VLowNxQ0WsW7WlG/3m6niufmzWmXZa5L8XFfe0V
6qQZsUKuey1Wpb9sfuNwv0yG4jenVCqydyK6pp7J6mfKGujA5d6BXU44IW2FGiVPmw4P6MZX610Q
AlbJLY8wJ4w0akhZ53XVEhEAX7qPgku+XtNx6ORQ6QkkGiKLj7tNbsOFqTM5K8VbyBLGmdfG2jNK
h/2lpJkauQAgMdG0Rrliqom1uSURvEGy2vSrNkVJ/69i6FsN+vNgi4M5yZMdbbRViEnbBMaYeG8b
a76Ry5SNAyj/+IxNUeg8p59xwNfO6NjTOBPIqlCzIox4CnUVelkSNfFGw3LTUAc49n25qCqvNPxg
NdTfXMaFhQS6ztqXcSDty0vsN3WpSm+t7Gbzqh8CsjKLPJUu3qDEE+VSi3RxPgKyB9LidFS799fM
wTq88y0D0PhSjR/Rs81y6gieFQJXx/kPx1vuQcTmE9jzU2IMIgfQGphz0xo9lETSzq/3fKVy1e/W
bOwDYsTM9j3rq55YrYSZf26lGJLAb/VmQ4SfEkp6+iaPfXZIqGrAP/M9IzJjw0QxApr5p0JQVXRd
pCp2uKBqWXJ20Pocdn+SsQzqli7hMxRR2QuEQ55OFSp2HIo1A7dNh+QVMo8rf08htNmelX3eNSEQ
K2eKo5PcPOkJBqYAFvUpBAqEn1syg52FKh6bBoEvGQdo8IRTZgc+czlxgDRI4rzh5nYaLOw6kHIO
PH9EMP2L+h9H329X1MfKjAJN82/PSWnaXZg/65lSlHKihBECZCYFznmN6xKUi2K1w8CXXZmjugT/
uVkWBdUp7viz9TP718ea5aAZqnP5rwt/aXxA3qjBD1qR0fZyYrwkbpFhdk6JxgI1ClSmgUdcuYnR
KkG1zY1RzB600OjUfwuMufO183swP+f5Cydw8kBklaopC5NfbteWYKUUPWp226w7uiFDOXtlSghL
Sa8FBLf1gdAFIh4+yzjLCDF/PeRsvE11sysPJys34FkiFgB74ta0IMfQ85CP4k+f8Etw4nthPdBM
mI7urLItgN9eJRFhXqLFwRl3hLZVZYQ2Gy8jNxnUkqEcW5NEb+1h3E4qDPXej+vOApa1wXrVQkpU
Mi4zDRBythLV44tuWN13FFI8bBfEBdrBdy/VPRNHNVy5oKfhy7/H7H27EEHgKGbZJ/xRa9oc7gSv
Igg8zRT8zEdMHxlTiyLKlKWT+tvolrOK38gxiFCATINf3e6QlwGLeQpZktjcAusib/92SGlqg9nA
o+o40+KB5WB7S+bk8bdqQCaOeMxIaklEPh+r6dtIEUWwCOdVbwDOjKDFV//xvurib5h6bA8Yp+5L
KYg/3TYm/j4x19vPiBTvhljHwVJ884pxaVgOZUW7wcYJ5pjQfGNk8OoJ2dPoXLt9rG05GvtSAKTU
w/oI90M1w9ghg199+6SPcSu7nr9YUXuRYxPwH1GDocz+6Ni88YAMu4bkiQlZsVhnlj+H7FM7812U
rKSOhdKpsO/BsPOvzh1WXbzhFvur8gXCOCSyCGnNrGILsFXL+23qTsVPKH8gUlOGlNKjKA4JDgLU
jN9+GXMcm7U0MlBGcSApB3u1r62qbc0v4y6XknC6/MDDN9fWyHknZ8qXVLhxig5QWd7Fj7VJvUID
K/APpyryiOjRDGcfvtdzHs7adx9Kyf16DTZREZEoqyGFUULNn/QTAdDdz/TC24nhP9ITFamLqDrA
Gl++dTTKhm/ZRgy0qVoi3SvzvdHydpkN0yVjGXA1krVG4e9sykb2dygnSc3OmfXAKvWrrsTKM5kH
dUHoAc6m6qoakk0rqJM8JacERzHb8JrT54MPWTJAn7wxWT6uYERoViYB5p6Vay8AaUEwKLbwZm/2
RCS/qtbhSje5c9QgHX3vlQR7lzktKzYGHmcMo+dO8f02RoNDB7gxdOf4DyoODYzZ40JPjoAcFVIj
f0za9y1sqy1MYBZYWkNQR5Li0bYbFFfRyVLScTJvUXJHc8JoQeK+qfTTz8expY6iAFwOuSlvfhXX
cTRG+WstBE8UhYUE2XQhk+2hrOjKak51kQzrCi5uz46h1ucaJwN0P3rKV3nzT/WfG99RI01kfo0/
UwdbyaYU3o3C99urZ5zjtNm76OshvEhhlkN6Nwjhor1kepBe8FtQcM08BOn8DBwb0RpBwgLFUepF
hn64FuFTian8mbzM08v1ePZOjU/oQ/u8vCMXXIgTmNM03UnW7OCBpzSexr6Pd6yQbCN7n+5HoYhe
h1QwSs/EX6B/gc8NAyUKw7j8XR6GuFBaFGK+oBdYurS5O+R56CldkD8p5GESyFXqZ0JMNPbJYHcM
QI9Ytk4be6RDRYvRNYFWn7F0EXpasm624Y+bU68EV2pFGGqiD6YEeXj+l+mRFayekNbnA5yg3iNo
anzgp2vmMHHWa1f9xUiapjV9+ApjnlMyE56XpiTL7WaGKHYSaGLU6iyLVkyqN7FePaDtefpYij7A
EJ1ate3BJlm8z67co94b6ICDm2efDdJOe3Ue7Zb4duTJpHubeGomhvf1fgpXdAFyLK/O/xD2/i8J
nZF3b6JK+q8zKDlofbJVIRvCJRwMy9RRzA3k51KoqjxduKZJ5mnf0KuxRd/KE2khXQRFz1fWXMnz
JmTGdN305lDNDjZ7TaI9/6egZkFsTpN3ZZswFqK+oECtxEKO19d/LDhSXXboH787xYT/GIGUQAlU
IfM88p4Ee7gzedneSicWxCgxwe8fFM14DJcKlnTn8mzkvHRfkZHXV2fO1fv835JrPBnGj0ZqYQbG
rP281trgg9oVWY8dYrD2Dp4XQV3deDIbbiWhneXUO+c8MIpI5RZIYKz44YNIhU0cKncgwIpKov/I
xoRds3grw6MRGpaR4Gs4l5mgzw3HNx6vyXTQPZfsN0/p0c+Wc53p1ZgnG8ZMFo+4oMGtAhjcelrH
+KMtwNrhFseXg95lI+yCV1GJdTRHreSWtEtbLUdFUux7pR1PyASZJ0Wgv93bhR7nHX/eAMX1Q305
eYv9l3O7TpVRq4hwR/fMNpreH1CiYlRcLi/6+q1UsGmPeUOYOsBn8FEd1E1NFY2ZojkFEg3pwcPn
2V2UK+/WHZWgXZyda/NtJP94jLL6wn2iFEMn+UWaGkxExwDqzvqff5nXQZhRPOIIs8N8+z+/x/gf
LOCCgnfa1eqT+1cfAzNNG9UBO4pNWe9LLFpn+dGn8vUEvEUB01TNkfai6xbbomn0m+gcDTe/5NNh
Djz1H1y038cPW8gOqy2DBqol+w6BvPFYnUuIEjm5Bf2iDoY5tKwhcc+7bs1Qn0sBxGrtfSfju9bY
CJLziyEvq2QjLRQYEdUaT6IgzKM9gXDBIGVhqmzlP9JsPZ2kX+OrNs1ySdo8UXKU7HCxQ6WhpF+i
PEBoTkMCqwr9hL0fG3G2YS1n6GuhivQ6a/GyXlCv4Tr6So5DebFcOjc1nwUrIdxVGt6Zwr85/P33
wzNN+WFQAdb4SZHApDTcUcTwdmjl7B0x21BUTmHX913ItgokWmwu/NoRs7zWOjqt1cRL7xsVAPos
LMWhqw/dsZFmjXBaMGpJctORf5v7g4SspQhlxM4+lFLOrraGHVDweyv7lFWa+R7bLe52h+aCrnBt
GWJni3jHftkjLFYBVYajZT/mynTluk+N+zZZZMH2TbBBDH16zfhq9Nk1/gR65qnZ6xwWW1KFKyFG
KBQ1V+9GMY+fNHLuqiz9nYkKL5smgVyfzjPmx3b4Oyq3mOTNgDqD8DDYymMtMWiT3Jd+2vsx9N0O
AX9kDVJTpl39x6nCXfWmvMRlo3yUvgGdzoiPGj6fLfsyaWYtlmI16zrKGJE6lhVEgzSTxn6sEe5M
5983GOoThA3EHXYJgZ+d1/Jej2nr65ehZIJHAcCZqYVDI2rMQlxZtR+/DTlD7ip7UMiUoc7mBbW8
EkOoLwokg2lxn+i3jXB1VYWMdhxwEguGZ4mxHd7ZnD6kG5UZnOCHXA/4eo04beaf2w5dmv+g8TVc
l4J0EA2mAR6+X8LHWRVlYYqrI6vch3mzBQ0EWzzGmUw6PsOruIcQA3AJOw8lctfspPursHT1b6OP
KvsGcoBNRyavrt60NtR6N3065n2oZRXEk+1dPZsbHGobZN6SSYkeD5vTyxc5jnOM7Gf6P49UXcf/
uIlDVINWrpxqtLjrcnyE7hZG1bviYJLSLwu15bqmrsW//QvxoF7uYeKYOk2kbuhgE36Z8PxPB3E+
fBhuf7sCIhMji4EkDSL1TtsAQY4T2cGuXORWQsnYlArYu+YaDoEDHz6uJVW9aJTJh1vY3T6wAXHM
bdZ7EEV0jLgMjIKo6yFEJQkiqlR9TTPLtmf+MHV6pn1tlEth8JeLLVd/9rUfCRueaGmlo2RuaIIX
v3p1W46MSru4LXkX6yjBbLp62xCdli1lbO2JBChrysfcXjUYezJXETr0WUJ7M6AkvF+vt8Ivqj8M
yZDqTo0gQcGSZoLgJZvmx3bTJL9lYx6MH+9HoI4sCIWncwlsEu02n5zO2WxJQFY/wvLSIi7x0p3U
YAU62sKhBr7pjNB4LhJbGp5YY3U6Zkrf48x0alRrRf0SwBJjaF7x9J3vDX57wTaUbj/zigfXMPht
dwQFb7d5JxRKPnSwAHiy8m7JXP7ocznXcLhx/JBqEJI0BBacKFPGHgqAxjQZDhwkx+ppzqXYm+7r
CUW00aESFo3mtxaoMGOs57y4n55/3VQPVJy2H4Kup3kgm5QawqqjT4/kzKmnIFvWzFcXzZEDYUzr
miETMW2YbkZ4U0dwCbiPJJ2Vvnuaef037P+vKasuhdv4YaAyaNnqMJodBHYwt5eK/i3pgHguY8qy
W4Vq+s0nXUCXsw5H/LO9HUP+6vVGN2Psg6+BaXQyAqv/CxLrBYpr02hRjIMq8eNU7kZJzdKDj4q/
tj3kLEKnWNj3I8KGW8WKY9zgsZaMqoVKj5CU1sQ82JCN1PG4r34B8I+0oq7BDSsYeUxuPzZdX1ic
T573psikVuJU1PNQbFilwoONV+Ri1Ie8QGg2Qd0cexe4vioZiw5DS07VfqBwIuiK/DjUq4sq3xrM
tgNEHb0O3PjIdJylIeBby9QpCvDNo1sgrgEbWqE0iSHZhhP/UeNyMTxWKbtgUPM4oEBuNbwG78hH
MW96gYjhHW1Ns5IIChS2lHCAiWR/occTQi4hoMTpC7J6y6vx/eWQ8UkS8ggd93t67Vk5vZeIHRHg
lzxnh1oviKgIMSv5lKGY8GyTM1IkU/efkL8jqwwuBk+xFr5QQImm/A3Ipo/Ur7HaumXUU8ZfmZbT
nlSYseQcbxy35iZaeVd4wNF3hF+p4rizag1ud+CHzECYQrPw8TUudSxkJypuIpKSZ36/GRSQDzpO
cj117uRN7Y2K6BH7pkgMG3GhN/qErDh2r4iEVa/nEDkFsReTIJigATJ9TO0CuLz6j0AG3HE/LPx/
ueqi562IOAPsQOXwfFL2IiQV3gPqUubAqz2sKll0VEQtLanttqacc8XBA1OtY1sOM4kI5oHReWfY
VFfW2TA806qLoxVJ0NWfg5qzp3RH0umgA6aYTyTthfUe1PUaMXZqsw9RaBfSKm+excvjcXncLwnA
a2mF+DZEwoVA6Pk7Z/NWGXf/ztmTqr3MWzR815273uAqaUxFqrSKXsS8jKtMmmfhc5U/f4tbXh1+
S/3cLp3UXT7THT6CDhMYPEZRO1B2DOamyo0pqsPdt48z26uO0WO+1onF+pGIMIZwUcKlRVTd8syv
ofjbvmrECfGekFGIyyELScgyz3wFq6vnVMI7In5Xkmblfnlm0bnLIdIKla7QkBQnrogz3W8XAev9
h1S5a1deDIXOqSjJxaXbe4GjIQjyZkzHgsohVnBza94VFKxhnZK5a06yDuVxuEkz8QkQA66Ff7vV
vU1c07PxOOgLMz+0+BMR8J37Fd4uZLy8Ox1jJf0JHgaXu6QadQ3P0tZjeUpwa1KntxrVouKAoq8s
9koTtwRUEHp5n+b8F16JJCiSK5V++40fpdugwqCFYWr7iWwTyodsyIEYj2Q/S0ZG69T9M9BkUkcg
sPBxk/JMzwcAPq4ydGFehal/a23IjL9qSTi1No/NX+wMWJyibvA3NZi40r/nnz+2/AuUwgAkKvit
j2V5ERQM17n6GESkrtmm5YxLljTBp83GBz6Y7MulVx/qj0okFrGniCHY95PL3ajsrSUmORSIHEui
ARxx3C4t7CL6ckqE39HwOH9/ZRuInd0D2v8aCatG9yVTQL7XJOqABTqOKKgdqZ8aNQxfENltYCIp
wx9K4v0/3P2NYKIt9kaiYN345uKd8YkdVNVUr28IyV1rcdlkNPgpNNUIy22HjihK1YUQUXwYAoXv
ZJAJ2F+hzYua9dxvevZq7tgXYpqFzYy7J3k4z31b8Jz/b9yyeA3juvzmgrAfhxxJneZ8ghU397T5
huLg/LwiC/ef6tdLIbW9afUNKihqX6ZpvthG5QHPPUOuIVCLhdiDA2IwT3Obf5nUAOFnSe9NJ5Eq
OupF5PTZthRRfKUueaWmfkFOkUFx/TtMUBCZc8N1PqKnBnOOsqEp3ibMcnUMKLtsxj9GUW9A3a/6
y023sozhkorU4AmgC5huueLaZcbvZjD/4DmFNcoqp93JlVuoB+A3Y/TXlHeA5HpRLnZ7MAuVSjuZ
+v3ZdyIzoldkdmq4Aq6oMAQPBp5miwYN6E1WALMAeIO9r3hnKJDvw91YkF2DOFYR9yu+QS4P+rgK
k/+vQStCnaQFt53nVu/PG/ErAiM7LouP43T3twLnYH4scQkki4k+bzbNFdhSOoVxoTdlXaGCXKHr
7wy0uBmzdywNu11zt/aaedmuF0xeSjrfoUVn+QYmBcuBnJfdP0oSelWTG1g/hmSvKOIkYRp7Zkke
aJzmDN9fVX7mA2JaEF+i/6hz/9cJxmqi4uLD18A02UoLR8nP/OEx1yDms0M3a1aCrypA4luJl371
gG21jh3QqypJzcvY+xaL/UkK/UOP/Ow/RAGrawGtSqFUPYTGqRBXKbrTYk/vgLh+0s6CDFrpZVCr
ILq+OQSbH6EILom7pjOaX3fizrMRHwl3khzXWLGycPW1ljmXOzFhSrkS+NFWuN/nPegRqqDcPp1Y
eukSZryt1RAVAR+HmqHfgcT0oCypiMGUkQbCLk7bksrpDyatJXYcPSOp5OK8oROniQAK5GovQfAV
0wNDC9v97c2ek2xQFrS+aZ4AK0yaic686O6KnH/iEp8Emvg821cxG6+9ExIFhcpvviodoOfinjCX
yimTssZjt0lFncJqsWCHYAMe+1976J0gL/nrfNww1be23Ir/C9iKBRA4bebnfH14A7dEICXAp8qZ
fpaJchGeNRP+Uvn17PhfOSxD6u99VZCNFV3WXEIPTn0PlmFwulzZ427pLQ32FhDwV9u9/4GZKZij
ycC9N7pB5fKd/EU+d+7CEiNGPRlo5P49qtvw92cLqzI8LRKUzSXGFQfXHZdAyoF/w+gFp4T8qb4H
HXSKSYtgk2R61a/rx8k2du0Av7+evJewpVhSLlkUkBdQlJAkVqbR9XqfHd+YggWJnlU5blYmB1Ux
Qoqx1Z+7oQc9wt+O5pqHDuljbISePh5emGyQk64r8eMDVbK4mVQeorC/SGjNgfDmg8fDKiZtLqJ4
CLkM8fC/Xdp2hPd3utXhh6W4mt5nhHxgyo7OeRbkBpiyAYEBrwtevxbOyZDxn8KPPuoZN51FAcd+
4wLp1/Adi/ITCcUIcmmEejicBfAmgqQ1jLNpJ2bsvB00v7WJHAc9pkOTHNsGzdPh79bJbA2vGtlw
yoKMPR0pP1cjso9t/wCYx0MYP2y9FBnJiPTVHCwNPSG6kQhq+T4VtMiel2YGXSyJ3zYZtpj3dOgz
wL6EB2DnhdblXbQ2txOqFROig9bHoq1WeNLiRqte6VE8EjKsz4tzRsrxZU8Gd9ef9zuXP8ST2mHI
NoGIe4wvZ6xghETK59+ByU4RWwDaA1Wj5ICpP4+Tc8zQ/Z/wCq3Ulj22s5MzLS0DqIrDgcsDTokn
7xssEXuHOg/bZ2v6/T2eNp7vrTvpOZA8j3WznNPMChywKSQG5Dw5bqHy+VmTivdMpp6CYTzhBq7a
ErkKZrR4TdXakjAsKpA0F3amdOSWrq/FNao4WM72Uv903ObrJ8ASlYQHRuje8w8HT0wGgjxt5E3E
ZHmBqJ4/9XcFcvVTd+s+peBwQSeWDgXNEyhDy2Ux4vtGhi/yBzrnuBy+wlEWA0Wsu5GZ3nSNzXB7
Fj7UYAHDmHEQY2MCh7X+2b3ze9As0qz2EjXp8riQBoh8b4ak9wwaqZzJK7zfd+I7cH4znFINHd+3
/lJwOpUVgqoQ2lNBYnB7L242DrkGLgMNn14vs1D2GvQu8yGQ5YvRfC6HpV1D8zZqK6+9fHuisZ0w
hkiaHXaaX896NIENua3u6AbcHCd6QzKBB4+NknJ1oulvlAgHmB7ijdWAwoDEslHXDdaThuM2/wwH
Ul/BxHTNcRCHep3VlG0dTRKZ6qnLJ8P1okgf5e6o1IYm1iuzfoakt2cgD/wI3JbMOemKL65jBBv2
5etFFL4tL6+CIO/zXUGU+S6sEv8qO/2CoKXUT6PqbFbFehQkofKQhXRGy+Hh1l5xEPVKBf4oc4ab
AqVmkfIspHJ0qawwzXpaCxIWgBRGZHEjlspsjhysfCeHzN3IDzKAkWAlIAjTue3ba7vIJlx9Ixu6
RfArZYSdzcwK++Lb1b3EVF0IhEvyHoamsAmWzB0kmItXERrrB8N4PUXSYLKxxEeZJTJXfMgcwS3q
tnyypKRhWU0hf5vSQ5QEOa5tn9Cba/kIgU1DcVbDP5XIjzWeBeM3spaM41Ub7Ngy9NTZY0dL8tZl
wPWYE6QM/zprP5Pw8gqoXGM/BHSgwpfQbriKOzj402+xl4fVpz3fl7/eaW4gaOCeVjOxN+H88UNa
K47KCuzW8E1RBwXYDH7EvvupFZt1kB29Rmgr1lwPgNC4CiG8COrblZfKxmRBj3tB8zTm1yt/O/1p
iG5XJMw4/iOxjT+ybcxQpiBZbJUThWBppc0ZXW+4uv7XgwB4fiLJQI9grB/y34zO5Ed6bICe0c4a
Br7A5lWhyPF3c+N01XiSv+/lM25RoAvcrw/q0uCQ25V4pi+MpqUtafBqnGNDiV0c+MJlKWDGdEyw
8l1DDcCm4N8AIo4NCAQNijNV8aWGARx7xi3+9quDjnV6MWIAx7DLR2rokbJTkQsGnAhIyihWagZ/
pmCboC+psWuW8DhPN3JFzY4NkfT4IGY5IZGee1IEWvhmYG0Bg72WdcnK75xo/Ht3dS79rrvLg4O1
XFxTon+oQwSJkL+9+m4kMtmtq6qBCntYQAh6HoQHZiupm94rO2HtqFCwBJiFn372rXQjfCp1GyLE
UH8sicU1VyCKGYQmv7ulC/W//5TWGJIDmPGZF8Vuv/jBp3tDPs99+Y6R7RsSByuB/navYNd6Emee
nZ7qvc7HicOYhTlB98IkAIOiuKJXBvCdv4v2A2Q8prTt4mlcepU56ICiTmRuPnTjZVUJotbgQeyU
VfRS6ZSltmzDt099nN9Aeq4CzLnQ4ry0/XURfm5Ha6jDdcXdCERlVyaBrXSYvxuottAcE5pN5478
g6iAMprDWirPAgWeZAE7KJhTgmGYHT9YUvzBjszBJ2uM52Oxb3MNjaHcFpZxbjkY8+vFwvV0CIDv
Mcw2h3jTmIw30CZ0LS9GEjn7O9/95W4AZ5kCyV1Pu3rwaQt2khgzHPA8xwon42dsamFW8cF2O8vb
LSHTahipiOpUf3jtXW9nMk4O8imCm9kg9LbGOELGa675mF+uLtG8PfU5niRAEQ/VzS6DhOAPXL4l
KOfM3TyTBhF3dcUuyDiasuBDom8wMm6wkqJWG4PFEggHRV9lAsgFYv644GIYu8IOmWPiDBNEm9nB
tkaTS25/w1iKCpWEko2TbYLodktzrP2fMTMFZ8irCXUcZ6i32RFj5rPDDfG87bIAdTf34Pk2GOAp
VgqZ1pDxXzAAg+D5W2AIE+TamNM2KEOEDJ0DTWGUyhETvES33tp602PD1TDwGzZZIEI8iDzXg3Tn
r4etx6uIO58YTaWap1tg735Em5JhQKj6cVXI/EVNo+T8ke/vimkleHdR0inc2NcOx7F3og+kFFhx
X8T7xq74nLjwnRav3SHzdpoHy/CnVrIHgGdmNTg7qy8cwBYZkiyBaEJMDcSul1KzGHxAgBMmt1yn
wOwbzBK0TOBql+yPiVaI/RcwBEeEzRwSTyxlcbk03G/zX9TfRUUwnXjcRr0x2SAm4cpXfH4YmwfK
fdOod8MC+peIHjMH98mviQqlLyAk9uFu8oEJOvaiFKEOdXOoPnf9oA3ykAWfqIyk2RIRfovOQTlP
0dzs8B+wn8fBKQnLF9MeKioJAADZ4EEL0LzbiDYAXrhgmEDB+8I8L2heXce7UaG3Gj3VO5mQGpRi
NvRptCzm+jblDniF7YT6w9j8fDS5nE9UwAVVGUtHBsDLR6IiqAPqCPbkIwUWNkeThE52rDqpDqD8
AaT9WhauLWwCW38Z9iWImx/D04HTIotcMGUE9JeqyMGk5kf5in12v72ut8b8bK7u58kL9nTgkfxo
v8zvxTvO9er/PykzrDIvoqRDX9Upt23DxZgXNt32kgILZndG2tMzCV9d7fG5XaVxhFa0XAxJgG2m
Z5WZX6Wp8+Chem2+DhxzCGK/qtcel8a03wvxYW2QV8nywnJRAaKTTqUb0Fx9m95Ttsz1nck0APBc
641fueohs5fQqocOFnhWa1JhyhvTQO1wdz/3vEOEttJZNh73z2bnrAM2r5VbHf4u2+PXtFmyfnzA
Y+TGUxBjTxcgg4X2JjW2glhENPxVKvFOCdZA7X0Gd9vTMvpWDVzkVFMN0r/QuxxDBMqKaxieVnCv
J8qnrXYoGJFyQBA0JXKjhsmA6h1M8eqSOGB95Q+Idhqr1AtFeKKalKSm7nki+TerFwSZ8t6elDeG
B4MsVTjzxpupleRUhvdHuB0gL36uEJ+SjO6JsmC6KYlV6+D3dCpC67/llM+Sbky/3NN+ye2YXhxq
stGT+Qmma0ET+f72W8y+z/4u/MXnSRYmt9JVGdNgN2iD7tR1S/d32fKMTaZii7F6uOWnCDzax8sm
RmB6iPf3buloRtBCa0CjZbYTzmEguQnjU9E925qOjUzcfdAZrX4mv/irhb1no/ROGJa91rBkBszw
HqNbNW76/jPWB1kroXEfjeF8ljaJzdknZe4WECV994CtqddXHw5FKv7PfUvxa3B2XA7NvOwaMAMw
yTaoEJDDLPHFNuxnArU21+JV3OaDCMjKA3gyppdbHYdipo5ARqYJPMCrOSx0zx+WIei9MN70UWTw
MApUeWkT0JpQGkOLa7L5aRxR7dMsfA3hcbYUf0eo9sE+5/SXL1ULx3HlQ1wXLcJBpcH7VhAVz00H
pkmkBDY3FJWD/yAin2qzLN9xs+NCyp/THEqwl1NocPrS6eVMZt/uuKEuUFbNs4Inz5bJ+RMYx56N
j12ZoMk0wTjKl69bPahc0D6QdztnTK5Gtz9D+ux1oJNWdxCB61HTKkK66MsgV4ea9VBDDK8o39yN
oPdTcwc8/OmIMeUexLYE81zZVDqnc7Hkq/Ep3KpOQvpIRYLb+HM5eTKzCS30gdADDGE+Rse9zUzg
Zv9lvyYQfiyp7rvWm078vjTFfYAKp/pVtUTUiBaSCP8LgfLBjF8gzYeUfSlBfG/tKJ7c9hjpYR3k
limrtqiFftswpr6y1dNcWeqJ9nZuOUyl1+iftQsFxs+krqgpO1Lug5QgXk8QQmTOMlVqlt0z//Og
kCxBTuDQ8qZgJJFQGhMlM/780BXUckiJhtgiI+gIVscgmUFLcv70V/ecSYIZOCnpYnj59gVnqbFz
Fjp3CYVjAHsKEx0IhzBD6K+JHy3jvhz7vazgwuj2MjmsL5hQtwkbpKHXv/xjdM4AF6aWEfdfJqb9
20DXNaAToz0UNbnz4JDdZn9wKVvskZfN0lCEZlvXZ0XYen9mjr/cmsjdZdxe/NrzMXS4Y5vVFwI1
DEOHVnymPQnYgM+vVAN1WY2RP3M+X7oGAansl5f9hT4JhbvmykOFyLal2Xa/pOJTac2L+5zKDtQj
RF5yC7FTZmEVuGTmqCKQlM0z0SSuAoKdgbJJ04gkFKp/yT3EGdFc6HdtImVMgC/ABSwVhPiWzOUn
uH2Hjr7sYTVHGu5U5In/Ykfsuw8S/tkieobUZJZxG9xJi7g3bIK2Uct+x8GuhFDVGNZwSndaGGHH
zyF/I3ShDl1Z9NY7sLTllQAw8ma3SeIkS5tLcPFXxOgCIQYvH19SnSRHirhy0G7drZA29imARCSX
ai09Emu/9SZ3d5QvsxTrTd6DV/Kz/XYGqNKrTxhDSSe74b3gtNwzB1fgs0S0BZH+XuzRn9Zq1a/x
mSdg/OaM/i8VDKPa5aiTicSpJJjGJLlIFHDujSWXwFWmVS+LeAeW5vVdjij7ogtWxKSfL8i5ES59
l29Yrf8ND7KND5r5NNlEDbhoS+j9MgbNWvZxoj6LwaMghfirKIA4PlDLNw3k+XyqDFnxhs3NiPHL
O7/BoGdIJDaxhECDOrBXmXm9sMKjccSdlaBrYEhonuCA2ojS5O6YwuL9o8EiekUdcW/odH+gGo5h
Nwa9V1HhCxJpyKZAtvPKmfhTprEkiznxp9cb41X6UB4wz6JRWhsA2riAf1lmhscm4PgRKsTLYThU
ZzQfs3ovrYCtAFuYnVBv8sOnK9oyJKRg0WM7r83SX03DxoVfXxBH4ID22TGLsOyvY0MY5wzTbmRV
WPaTop+eTjTU4jGJq3VtLPnBf/5w1LIGpMQEdp4o/v9YzFf+eMzdvl/U9jQMWfki7uBDVSJ7eKIp
gj2bwfIPsBy7TwWWYPFHL2vIpJhF1fBeXEzEpEmAQ+a/Q/hT1gFWmgGKl4f7eDj0tWlhcLEljpA4
Mjqic8b4R7DkeTyxt9XytqxtM8rMHEHuJ5KLVAN09C2S6dsLeGtQgo0GDbTq0oL+nnOf3dVYBQvY
QKbU6BaC7e6rad6Fgki9q/T5TxwxF5iuObrNfON2qZaSPcDZLbF3JiU7JSyG6dy+QzyAsu0N96KL
uklOUJf9eD7IQdKURwCkDovZjwR68DZX+24U7169ojMLJKO2BXUMeJj8O0Ev1+SDyg9EiKIA4yzi
URPlMIaQyeZbAazQjXl/wlqYo+vxPDBL2txe2ekEsU3ecZHFjh9yZ/BB+zry/QsVpxUm+iTkpCgD
6RKCarOzkkZZpyT0l/9B7bcbdDh3BXaJQv1/kVId5jiMXgBAZbxgH357yaDuQQjaGsEq/iV1eLpJ
ZNie6zrV/H7sYapFz9zt9hdtki+AX4OWn9xwncOQa84PYoO/xu6Pk3KjWDV4ZA972GEFomxoCKGq
0yd0Vrsjy/wx4HQlNz6l5K3lpZh/h1sYC1tpau2jrlEI7otEKcZVz9zH24yW4OBgta+W95xgA87L
waxKPrGc3EY+a9UfjvUnz68oqA3p3mrll6bOb50/1RnDaFKQsyLGO9xjeGCsULhiwCunDn9kIQPa
itq1BPKF/yDrDhF2BkHf4vdYsg/qFMeha0UWX9nt9ZeSngguwPwkl8M8OmLvcwdYUiIKfeKBWf6V
I3lQPdEgDdYjujZbcpC4LaIa4lZL9GfT52sP7mQM8GPoRYrLNMRbCTHM7FjF/9KHwkOse6tMf5Hx
w8qlH3DrXc9m10gRH+3oXlRvAJE4i8ovwK6sdp87T9tJFAHuhLb6Fb0naQvD0lSL20fNf2oAVbQ3
RlTYiiF5Vqjp4Il4x58T9HNQjvSzPwcFCGK1SspPA0lcar8bdhaqsLPxDY4J7C6Y9+s5OVDQOkE8
PWSQ+fA7TmiEadjHj62BGCjWTwMLt6gLC2zVOoM66w4/Fz/41nRKcIaJS8NeZgFxVr5VwMfyB1v9
4IO2Q9YlBTZ6Vl6GnKVj8e/M/k2H237X4oDTH1gBNw3n6Rh1QtqQWmZ1CUog3mNMQBMYtvYNHEFt
XesGfUBRSItMB5ItPqmSZy5GRaQteSrRa5MFLW8xHBQFkrPk/cyyqca7OoS6AhDMvcCbKAHvG8SL
58G8n/sUiEVEOODrQgceuPlnPMMr5l1ezR2A6X7SbzV7mTXEYhAWWHqAJE/L+h6GlyDhGVS+sXxs
dli/gnvpybFCDA+VYantgA7ucQLPuxwLEmvseEKeyVSVvkUdSgSo5PuivzUi4lnryQK7H3qx6UNI
0jgx8I3kIeoaRPqxFKOl1Q4N0ReX/xLPgfL812gS04Hu99S4o4F8elfdRP/dv5lOOmkq9JSOZpq5
JiNHC5Q4bnF7odpnHZbHcdiCQeyapKQR0t+EgyzEGpuBBiYRP83KHay3/eZoubtBqYZEP+Vn9g9d
QYdrJLgSA04hAPkfO+refZYalNsjdm988f1h6dl1mznak4EvO0JTmzjwWC3GrHba/XOIutq1LbhP
ZEPcYpCfuok49iUwbETJGkDsjeUF6OznGwx2kwkg7Yj9yM3g9TvMLWsrmaBa2iJKqcsQ53SQynHl
qN0b3Y8PH1OJNhtMTyDBA31fP4V3iYniHpb8WbuWX/q8iJoyMLZzfLY9ECm+e+Kx1lNnyjz5QI04
t1GVlo9CWObrG2XtR9GLmPyCx5HvOGNL01XaDc1DyNbxM3pi/VZB+PB9JvI0POz9PFF7H5S5wwLe
J0+vV28EOEXMNz44fe+jRG4fSEn/uLIC+iubGhT2GruIKwln6VbHOYcUfNK9eVS8xuwDmMtseVbA
MxK8fOFnAWKb2jNhw8kuU8aVx2O1KI4XNtgG0ymmtOEPs6n7BsXoSzPJTWKBB4LXwKoc/Kq0iQmC
9oYbdb1wpE8faSauS4cleorYolxdVl+3wsDgkpMXdlBr7Uq5r15wu9x1kGx8JLY2vqsvA4uQvKvg
jFj2U9Ez898C9EzCOyGU6+8qTWWcNCoSTv4FkruKxEETdFEN7214ylrUP5rQpPPa948ep4h7svPx
EnxvPvLyg7ISXOkg5pwLH8ozGdOx7SO8B+jPGNnwB4LtKSskcqbFV0ZMdVQOT1NtYc7YuiSmn/vN
MX0+lLoS5syTkxgwi57LMtyCUNbaCAmX5u65X35Ps5LQYZp7EtgwADy+eyKbpMi5nTDV8KWY61Sl
4LwFx9DJlgndLVCjVruKS/mS4T8D6UF8tufhQqZDjmc/YdITrBDfAVtHRSj/OHRk6a8AA4kBY+16
B1xyE+Hr4YfDj1K7tbz4u9nGoZcDBZBvekBN6ZmF0kxTUaezeCiKKeBpiFGHXbgWkJYiA5W/ribh
ugK10t3qY8X7tBdUja7koRSQLZHVakWPL9NqZzzVyF/v+scNutMqXv7uUfatlWixRsxdywXRjZVd
xmW3GENAz6JIw28tN+uLxp8uAYLnJlrh+xJCE76ECELMrzNbwFEds43oZnQsp1jYO3DVgeM/XBiM
SU/YTZJMrFUfRLxbfbfpPNTSRu0UkyfPxxPmQkdbBwJmrjju6dMX2Jh4eWpPYdGWAvOFgEcqkXhS
84bRgLvdzTxPuJPpY/D8AypBl4zoWZWIDtx3UoJZTuAnnSCgxg4C0pyKBcgxOND6ZMBrkGfiMIP1
wY7WH5jG/ESukschrQbpjG8Z4ic3GJUNWfPUj4L7oGywsrikLZfgm0jM8Ij3eI73E+9oRhBtG53s
UIPn6/1cTz63GYJWyEXJIJ03RX1CHZEn/AFqouIEwZto/vjZvKm/5ME5fv5KE2rI9GD46BYDbfvC
TkbQuec1Tkwlp5/wLVDJyMPSr1Y4zt8Nze5Vh8i28VT9jjnXdXD1Kt6OcDw1GwQY7LkOQukcYUL5
ujWSAgKCgC8tSa+CJ6yzC2ilplwlXEqgCIt6AAo/Uvsrt1x/AQLEXxn/ruqv/WggQZbi4d0Y02hb
2YS6F8wpgAKiMUNqrmZ/2TocYc1H/SzrbFcU7gXaTEDECkZ0Eh3r/PexpEzf5Pmhg4fKopl8HwsF
QFNw2+BbhWhgzBZP5VpPtNw0ZfkTq2W84ooVqDMQ9BbtOkWvpZtBE1JTXMKVUj7Jj09TRqtrXRFS
2r8iZqEHPDyqWvxVGKSW5aUyuHE9vLgpxn3B9Oh/Nj4w0ndLfoCmcU3iPGNpkyKPMTAntAuYvy3f
x4tTcmyAzUDaya3+xyHQVBl+wkliQtkhPRiUt9PC24eCUZ3dCgz74iAOdrUHQaEKzv8977dgry9q
ZX+ZDvvf6jpouNdO4nCFEzjhnF2tNXZFwL0MJ/OA4QdzejPrAP+W+oyBfE7GJXF3I+nljLs8IND8
nbHqs4S7afcaLFonzDi8xEk8knvNNT6DluOt2pfPqyNJt2+lgVCDlm4jH0ykS2dRjgDuBWGYooz6
l+mEspjBwoQMBeQWMVyHTrBpl1R4pRi/3lDOM6V4/ZlViQ/pkKE4mFUS8Ed3HcqGWuLuCbRDyUzK
q7JDn2UDGKaE0jbdf3S9vlS1aLXWNtAOy4KDEOwYX/eKOnaYHvj5+mI7OGuo6hH6TsAkgyX/u01H
uAusb9IVbyqd/XBDjZU8KuUU4M4pz/4f2hHuVhG/AbkNvsIo3Woh0y+ni+fymGWWopPBA+zf0dmu
Egm/slbZtTMKjrKDemDaVosFCrBQi54/cHigR39Win9z/4aa+RS6NLKQULM01TIVu96qSDILOm8B
UoOkhNMVFZ6H/05NWG8FSB6Io+TdDd8U2uL+wqJOUERICvVnnY0TRLZNOaEJ1vx5cMp17QP+AeAA
4CqhaRA4jvf1hqQzqgI3F9374BvbT1+qI3VtktrFlBmAwrj9/BJ5bTn2z8LLzh6jQQKRrJbuNdsB
o0UfrMHxgZgVozQnwK1GOLkhVITWC5BUwUsi52RpvLZx1uJOB70sPOS4ypX1d+3ZOG5mRt5sfc9M
JQQ2SA2/vpguvUr1L1wHaYqr7JdVXR16Yzuqsr9mjMwQ1lU8bUDcCawIVKxCMUc+25oJznhtBZPz
ROgLL8X8YdSOTsKKJE9FzonVQI7gz0rG8LuFHURgQOhYYd8aDtoh14/TCu8MJM9boy4UbVcdvcxm
QVjeI69CF4rJVgmWCkKGGIsVsrMNYad4LJmqYFFWA/q0tYl+1puldKRN/IsMruaXyQmmCKGd+Yip
5vRKvYkwF0nLZUp8q+MLCH0cK+twYtMyLntOz7/Wp9G3yXN72nFdpD0FX7c3Ee0bGKKVIxNO/jhu
1T6cWEKoc7oQkQgjairykEAk96dDgPlVOaWEIZcG8p5LicqbOE0k5mQ7CVVWwJXIWyWxBOTQjy1k
u9/8lVsrmQyjwZB1x/1Kqf4WJrOVaHHP0ekfb6YeV7CMU3qvoUeuV4UwPhifBOdUrF0ZTateBvT1
3fol7guxhY4R42SmETr6qNA0iFucJvTs4Dv9n7+m3OJBAp1QI28OPvRmj+rK0AR8i4qrGd42RvG0
OOF62aQmtvbW5VE1wfKpd0upinzkLYjuIU9LSVXY0IGofgitWAoQSF42i5wzPAc6jy+UB8AmHZVC
wh6iJXRdHVnCfC1eAkf/r/JV+s6B7ovmw3ytjXJgYr7Mcoyr14nzsc5RukJrSLidBVsRupBqtaKO
3WPDz5UmsLqn6iWlckIBt43cX2+CcfBNUgYESK91+L7Owt8rOS+eCXJXttWBr7//zzcdl5uryZbp
g9DDx6qNW0ZA+LUYTZ0DZAQZLiKNbpTkEcZ6YMny6XoEi5KTjM8OlGASTv+q3Jxihbx8fhUs9OeJ
nCV6qw6ds5wh9s0UudU2O/O5M5jHH3iiT9bKHZi+4n64jkb9HkWQQlGAtxmxeyuYrea1iCgFQy7n
tVFePWjJXlwExKnPNi7R54TNp+j8xEhcA0z3BQ8L2we961qhDOHDxJFGkMZCZzSuOY7wrVcuTAi1
yNRYHGu/TF38FxP4mP09GgiCQHB1UqCz1Qck9G22FKnkCcvEhaxEV2xBV/xO8AvaVcUTCui9b0zf
F4aX56PorXXy56ox+lLXRHFFvP1hj4qYmLLqJXw8ZCABCsKQxYf9HHI6rkzX0cq2+K6RfS8wHQyT
HBH02x1+m3CQG0Ay3cvyLkuQiok1Odk62wyLFSd/i5XOztTJPRR1naVPHUFDb98sIiyh2T/DFvju
SHcKsvnQYcM0rPJ1k6z/p7TcdLe4MJnqvi1umLtQi1RY8ZE06pOzCKfC09Eo/E6NOFR5zOUdPhqJ
9eZrAxZKcBBqBBen4PeKTJOvif4myvElkQ6XSgYK1MtzbpR8pxI9MnTzMZXY/4djP1eVkZkhM9dF
CQrrQPhEYbS03yXYUkJYhXMuzfClwDr/md57PESA4hd3h76rrOOiodnKobTxCX6hwIl7KkFJux/Z
VGaR6C9WMYVuuQNXOJQ6oifKHDjNFflCJRospbQZx6dO5gsBJhBjqezyzD/50PUjRt+SjnITTaSd
Cy3SPr6If4nBFemhzDDdyEyc5hH7/0e2YzKMBmdDgQcsJeMucucnPEmkwXB3TNsAN/ZZU4Kxvtdm
m8mpMiv9fK0hFIdbY6nRs0iyGJnSbiZZN4SMyt7qVLLUOlUyRkNI+69c1jD16nCjAsGi4KN+DWhY
fLV78ZEKnDZl1RBkYw7l3vmVdQBxbq4j+xaSL1zNVi2Aiy5e4aMyqrMPYTYmKfHJZgRXrGhwbz6r
9WWvGVwNMd377s8wD1BfcWl+xSKLiwrci7sdiPzz8L3gElnHBoLgd3qPsIwgS2qv99RemyBBBhZV
nnXv7jH25ODpnLQWoAvo8tKffoHuSBk2YNFeV6PoZaL8on/BiGAGyJC3IMqmrS2uG1Y8bwnqmUIl
L4cy0F/MJNHonueRjlrBXJIP0ADGljlewyfLKcIv32QKg7jLXfhMx6C748HlTREtXUHPQFuYhvog
zUIcTpQocH7XTDrjzi/wA+olvGM3XMIE/zLZ6Q0z6clohyb1dzISsmxsCrdYR+QNDUCC/uNySwU3
ZOVu350E4XezjawDxwmU3AD6aoedsb2JjWwEVlhP6iATsFNeBlXxPIYkay+4rSG/D0/aSniO+OxR
HqWjVCJRe+WLQ3YsJ7slymVFUR4Jcqhaw9TyYnqgQGadS8EVIe7qDQcRJqFEHtZE7IZvA637B9XM
paBXjqQggUUqhR8zo3wAa2DO1ipMal1OTxMYoYT8wEm+yLK925pxUPywx/i7sioBRJQLqqtIQFyF
jQy/RIZyIbpvv2+Dwr744LNfsza2GRwa9I2cU9Xl0FsNbGZ4EnkNSw47FbH7cpGvhXyDPuFg4PGY
RuHQFfz5YplBa+D9z1PHNmM/7mTMd/AiShgzC9eGMOVu9eGW5jqcDwIJyFtJHd2zHpbAjj3NS2BR
jj3mwaoWNG0LWuQMELXzRVuighRRJy8E4I5SBYduWLPkCOig/J5o98I+iHPA6l4QV6GBdWm9nrUW
ea+BapTxsEpc0pxFSRdYEky1enrHFCY6uwV2/opT09pS92cc3o750Z9f0UTWFPzMgHRFTh4XBVYK
+6KqevPzdz95Yw0EWYjas2qSYWnzWZnHXBkReSPoYko6vrhpPU008L98CMJ0/xQ4FlxeBNakCdf7
Bcl9Von38tAO3dznx5sQFobaSR+8hq6rSXPjk2UsdHuhsj1sBl8+7tnrM84LOMJVIDsfrjagV/DR
U19t2d6PxrTeycM2xshqogdLeK0sNymP85vmdz3ZTVZgwQ79Ta/4gjnHHrY3FAqdT0y4Cop0sLTP
PZOA5l/1qyWO+AXFUiFhfckzddhYUdoSRM5QJ6K2GQ6/DFtCV9Cx6KAaL9g04YxNjpjrIvQpmYlE
sXO2kTLEVV/sxkKDlm/UBfvZLuCU4+pLsDJjZhgoGWva/3mLHG5jb1GrEYxe6dEAOoCshfDMlap8
zpFK6v64FQmPwoFMfIsKEM7QhoMHaxgtcqqdF7MfR5yl83YZLgJLuah+CR+YAy2WE96PAU0MDXBQ
b87hc2GquWTAG+yc8z5TmeTq/UHEFq/aPoEeYDPwTCe/3uq6lILexLpPspfRV+FWj0WjwqaLXTu+
umkbNEmF4ZjyznmbJjy/UjJw2doQf3COU5DypGSdsHOkx/6KUnMFa3WU/MWBNQ9yGj60WSgx+xXP
lbdz2KZnkxcLIvBS96oywlGoSQ7z7mvkiPqUj+Uish1iFu2To9ZGciWXukJ/iZgK1rGcU81owbCh
B91kYwhK5qgpw8ZKkzuqoaMBDMW/F780KjA9pU8adq0sxbNuo2ofPbYGa939128BvsrBqA9SkWBp
1BSkcv5/P76dEVRe4juFkzme4Aba3CKK1cobTnVgtfilSi0CeEAZaaElVJf9mpNqNzbYrWqtkJCf
zef2bce1nlnooMDb7xWpT7yKY0+758j9A/aasZ4j9W2oYRE+rWkdaVq98+y753/K3IaxyihbSyP7
RFDqz8Wy9TKvmSM9/rTIIBqoP40/BFdW8nhVlHEoT9rCzG9MzSropBmrPcTBLHVG4TpyBV5JSVjQ
is/5SG5aFkwgkkfMmxrrfBxPe6hIS8ppKySZZ44A2hQXTMMPGR/KLqMFEGiGJOOvf+jmnPYlnANQ
5Ye1i7zLF1wloGwHw16zM49wMk98D9WlUBstV4a6RFBQPTGVrwPE6woXqQ6DUKKnCsfCChwJgTqP
q1ShqOeoO6aVyJMBiWhLwtIxffP4g2J1n90fA+RvVpzh84fCmvOu+DzewU/I1mdiG4a3BX3WP5l/
oMOZIApV0/2aJ5oB40xnUrQZiD+twsofPYlym1nrWo+jsFTY8H1rgk0YR5/pdWV+19jZQcObbtR9
vsJcit2Z9i2HE3CgSRdAK9HABmI2KUprrgTCjBz9gRbeJS8iwmUpnkMXYtWonL0VLJq/42NXC3t1
AZ9ml7qVY3L9ig5TPk6sbJid6pWQot/GPYVxBvAQAjDiV46xih+XjWOu+4hIs8pMHw1D3XHNaBbF
RVC+2nLadAOKJJ9lAANZUHa093nbSHt6LiGouo4tPq94t/+ewDCQs9PSiuacoVvQknv7yH+IbRlt
Sg2MrAiUAmgN3HAOVcz7kdxHL0QqWT2o2x5Z3vbMC0eAyCkRFoO+iKygL4oYPgVsLF67MjEn0TiT
yz26xdR2PSLqY04vMPvyvQwfhcodhSBowYqBzzDUz++DJV6/rR5EkI1oagUHkW95l+447DIqKG/5
MGTGlDaJsQOW6LA/QN1ZT39SfwgoGbe8yQGzuBCbbLNHJcu3SEDHpBuUN9y+tmpXr6ZmnR5hzbPT
XGdsJ3JWOzpeSSV+4Kp2wk+xdimhpl3J6KJKTdVai4nXz+zuIqSUMBe15h1TwgkH2U4PqtnLbEsd
TJVMcZePX6M3DJYNvt2dhPi1GTXM8I/mGgHtIEMEAGw6r8GHildfpqJ++HJ92zFTvSFtaFV1WCZu
YUEha1JhVZnDzsduuRpEWMJE08tOMAtPTEihQ6t0IRhAtbCRTvSgkvbjgraGYI3pd3BLINztRWE7
okFXp7QpkCNFcgorLpUhjyPtVRCqlypQl4DK+u3RWl1dK53o/AJ10ZC5jjYcDJ4BpIMme5qIK9HR
Ps3eXKuZZf/eregplfMWNb4hHvrvpG+iPG0/1LY7JF5DqL2+jLDhSLq+S/PfFleDPl6iJft69v+p
UbPHDSINrcDxuch5kCQtkZyUmum4bmfp9CQ2OtSILXm07y/tUOm2+I3hZOZyqGD/BOvHgBTGXNNI
m0tdde7bOAYGL6kYcFISF6JD2bQ1IHB9H9/083iSpZTCkTZMYgrMXadAxbzfH364xRDRLFp2lwTX
NzX0AcIis5LDQFbYtQ/yZLwkoakAhc8fN2rJ8SwU857ZfQyJks23EA9CmYwQPX+YQYV92HuAkRjO
2aUmP0arRJnzyBKbVV163RoDV0zZOp4geROFUc4Od6S0oeg6GjOly5NskSVkQpYi+4YO0+sIdd0E
8OxAWq1n0zkRB2KhYQD4V4KsOQOL7Ny0kc5k3V1kqvVFT6yMuWe64oCa/KBZn+MLDAIv/W+1041F
uAQgh3Jce+CIpc6VkQu0h5/+R9LHKD2XKDilFRViXRel3t+qLZbIthFuXntjPsWHHFWoHXlm9tGG
LtlEBwR8EF1njBpbPKi6LfKdul5KjiGI6e247l67YmDCok+Y/L7SZ0BlNn9L2WFiM/geuHLAUrwL
7Fu2iQvnfPIVh8Fl1mv9WQ5AP3CWpVG1bbl3P3mk/99vKEq4jFzuBUdppzbhz4B4YO76O/VHdNrs
XYxF52HtRaPNZV47S2vwGAQanOEOLi5itxmMWxDV24nwTsur/ic+GQeosqGz+vxgy5EATyO+G2Xb
LuggfuFga8Bk/b0cKBBOVjh3hwRzVPHM2iDNnB1No1pcbPBppmk/pWYd6/5+5AEPG/bYJj0cwEaq
vo9wrwL8njViIF1EMuYcTynBtux6+d9vu+eEPJTi69ptR/ngMuSQu3XkHCHrYSRex+LB6kyfkgvu
3GETuYj3h+YLwW5GtSjCCZPkBLcVZmmO2JeCZ5YpSPJek4tkY8S25XG4ZEZg0SfS7XFO3egx5iKO
/j1fRviktxBov4+lWW47T4UQFLrOFQEDFe7Akj63V6/dcTknOi5puB59V5MpaYZz+oUTjYG4lnkk
Nv+aYmQKghFyRbR/akTwiglOCGo5PAC91kvGrN2WltKYFxW+XP41h6oWO/qrxV2RWVbRnPgOqvXT
DEJ/fo7jNKZ58pR6g9VyGfi61V3XatttmtKuJ61jZZA3VfdqouRhSx2y7LI6AmsOyGDco7cP/3d4
RLfN/C2Yp8+na49Q/EXr6tvVrM3+6of4bCE0LqAv11NHiTrqz0Sf6L2dYUm7g6cM5gICV91r0/zS
y4IU0fgDuM+U6w2lDJdKV9pg/UGtrf4YiXAyRMwy2d4ywhLTki5WAapKmIwke3kjyYYMBRFH3IPK
kAyfg8evA8d2eZvelasb8AAhXiYhEd3XM05pX/SVbQYI4Qj2FB286x4OEeWX/K3aBKgKwUiHx/s+
s1QVzni5dVMy670xWOkCV8HIiIijLAQy6Rah6nXDg0ZjKGL+zaS6q1veOIkIWSi+KSlrKiqo5tEU
cXYvJwD4vMvM6wUvgpkcToCUgDGYcVf0R1GJb7pCRYuI1ZG9ReGCh6GNO2Du+SS/UHLoiRziJdHs
eJdrY4lFnGkXcWd3XAxZJijPZb08XGbUEzxBAQAGXnPiF9sW5wc62yFNVNBkWd6NmCWXfwTESHqv
oS2IQvR/QxraRSV6EO+DdmkITLQN2EPLRo7A/aCFyPp/wx9Aa6ngvDIDoiWxa9sTrLl45LlFXdq/
/B/SBe5of2Y7IemyT5LPnXHvt03Z1MJDlCE8++Cp+Pb8ohFViIu47GYS4k5gTMNn2WJT9Gcnruf+
SRY6w81lxMh4fyyV0lZU55VQDwtpY25tBBXANImnNkNxGgc7vWRAEYBeqMJY1QENrwb66Yh2Qw4X
yz+JvI6t2fnXDSuKy6jPOpJ9GeWzlZKPuABo0HiOz+4CY34v21aH5fKOzYyq94zG2V4E1Gzz4BO/
QKEyhCs3p7F+plQcnAh4sMvQOeFdR3BVVU3dQXkLCn+Et9Cpi5paFKwo+PxfGzTkVclQDMjBRd7Q
03BA8THOyMM1ROiN7bxuGhJliNtVubO15Jjp91SWtouIpPgF/G/7q19cJyB2noA+a7UzgRruacgb
ZFu4MqwJN9SdBg7oovqC8ui3FxnSQHGEMTwy2gyFzhoJMvv6OsuU6LZOvmLcI88SdHzbyO8PRTsk
wy5+r+djgCvCQ9AKmgp+YGKHEATxcNzY4XXxUmFH+e/UjJcjq1z0saL/uPzX42Wp6+wk9qj2LpiG
uzKyAH5tdKYYM0JyvYOzVH075suwND1T8tQ1kwPVVV9OJvJBpx9ADL8gHI1sTDT9SlnW35sajudg
wOhcPTQcEHDw53GLq7JoJeXxt/MvoRfIuDyU6msozWUFRiIHfOjOqiXrUIJY0ptdLsupkzvM+Orr
aD80XbvSKBDP3Z33w0A0MXcH+1h7b6FtpJ+AenBjERaVGiQsaWI/+CklOdYcHHrlCJO+KvW/K8Rc
rMWcgnOYgs2DPUTbV4Y78xyWBaS6osZ4bFjdAqmhBwzM0TrIb2XrJohynx2gH/a6cX0+UVh+EP7S
FYIt7PVXO55NrcaUWbmYqGzZ9qI/t8SwTTI7/rLnREWoBfNkV8CuIy9dVVx/q5+kSrwh5aWV58cR
GiuCRwOOH01SxYLgVcsUoVDA1DQ0Ra8ipQov1E+olzGafTl1XoZ+ubn/NsG+Ur6NCwsbpHOuljFM
AYvwxVJKVhc4QqjNvFAZN/yqSuIf5jNXZTiYH3ySuLPdZ+MGCUmvF4YbaQ53FHk56MQ1n+dPgRHi
NALJSgazhTI+VHtu5LvPxeM8EmGHFr4VYGSIGRujnUCY7K7+awvlJX9AGCFW0oa54/0/N8gdhOn5
leUKjig4DGzpZo8nQwmA2QTcG0VIU2IUSkxY7K7lgLX4lBzQ45r7Pezw0QFk0z83FEv6lACHKfOr
3wsss2MHhECnnrdgM4oeoCXWVtsGPBDD8r6M+pIKcunonmu38UHkaATFfxWogQZc2ybBdz8Axws4
I9wV+lmh3OleO2e8yeHR1df6v9BthStyqr0VdInWZOLVG6cslwOpj0AfYPcROJR/DvuW10ZufNha
V8xyat5Bhrv7LdAc8nN9xc+970c4oUgChsPUn8RInmTNAF6c89gxD7dpLDaXmjwEBZMAQdDHPId+
KyK28xmV235EjiuVgcKHsxEUeH3ibl4vStLUBs1HCUe18bZvYl8GSiCK6tCd3BV7CikkDAX+aUG0
wJmpe9OTp/oqEr/t77lllo/I+e907zMms5CSLDBCXfzLEU6+tEYxurcmEOWliHEnjhqHGZc+jLki
/V6f/YR0LL/3nQS3UNh3M8vpHt3GpN0Xt/QXNU/pieB132SiO1HckSBcr7GFN+dlRh7Q5+cNtJEx
xRBC+94dMoBL8PRly/6YdOGpISLtog/2jUnrJzSMLqxtW9k6h0supCB3hD4NLSlYuTV4pdAFO2Sz
oBxZpEh6hS95yo4mi38QDkRsuAykwLi3zzRIMvjloNSKt0IN/I0z503vgy2/fdQ71gChEYVXJK5h
xxCaUqmRiLm0M549EHEvqqRpr9DlBgCX93klH0HBo17KIr1CqO7VdeJGleL0aN/i8TGqoiERCcme
TVgc4decs7I2xGH9BurfUTLhCNzhyyXOwk/Lxz3/ZXA2seaW6NPXBUAQGMr5esNS5W2Vtw8u/39Q
JYlHAUkoiWBqWJWbje78O24hja3ukSZUfXunx3+FR8AtLi1zLiQwR9WYylTMGQr2RUZ7sS2g+6QZ
8Pe3WhT0PcwtOpXS9HtAQt4Z9y7tA5tBKTisueqPdScllKCNVc4U0OJcFU/GKt1ZadMij/xGw9tb
NZp5/plUf5d9Vm3vPp9VfkaKVagUf0p2IQlzXPmRRY7gPZqWnvJQy8DYUh+fI/4KI3sJkcE8BJCa
TTGNdKctiWwLVxQNDXBY++f+twRW//uGXU3uz8VQKNsvnz+i+/tOtDupBM1O8v+2ivbl9XV2OkqP
DLHJTr/gCRsMjdOB30prF3gdaqUOAg9i93/am7K4+q6VnWerBjigSoA5naVjDF355NbFBrodNrye
NIcfBbBb4BYeVTAkxoUbyTQ3SkWJSjVTy2XEGSkgSGGJTfpt6+I9no7HWNAonjlcjZ9sKSE7PVMR
qTHVagUvrDH5RYBmDrDhdj2KVpE908bxFJBRaIONput4bHy3y8Fp6RHqUYUE718PSu8tdelFglAH
JfJbo6wCyIzOifUOLTzpHPIekrmVQF/Wwh83Ot5e05jn3Q0EjXYXhcqoCPlzdMOzvz5HrG4rDAaU
6/cFEbKunvfw8uYAKn6x5mP5JaVp4Lbkrfh1btM2eeA3UBbAchqY4rAbhUZZ28U1NgT3q/ldVtJs
toP8LmRd+h444970tM2lBPvjGC3I4Xhgn5xksKN8HtHAeD1igrzTVGi47+Ei8c/ymNn7mXAgV7wO
UM8z0aJY5N7WVCgS0Hc8SUUboLnWeyDlk4nkBfMsZyXPuR/DCKZzehCOdzrOn2ohzoDBtuceDMT5
eAA0M1c+rKpmhcikEzOd1Od3MhUR9uWNWNA8KTukj36mXyqf4OykDEPG1RrElVHk2na0tenvgfXA
FTk0NUBsmCGJxlb2i8pHngWMd+wfuoSUz+7aqzpvCoLLhm9+LpQa0lQHCtgdkIuJeZudpvX2luiv
/xOhWLTTpkP5GHbsnJJ77mx4mzEJVVeR+t3oD7BrFhUpeqI1lajZ4bccDwxZ4g3D6wk6joTGCBT1
PFnQvPCL7STuXnJUZqVxoa0OMtgmk8Eeh/DQ9R5eNCd+yzAeGAnldUlNQxkHKbqCkAp5TmqWdWXe
IP8jHB/c4vLCnSJPPJunz7DIEw+uSeLeH9HHFbCPaUvpfklfHDvCf8CoszRVsuxregDlx+VHIp74
z7uFuHmazgaaw4GFTa0zwCeswQ87CUhGhF7PJ97Ut6Xy1e3xkfgj3zJj5yD1cOzyvEA8qQEAymKS
CRoB2fO/NgHup3HdPixFODowuCPrH519xlOupj1bc6D6c3Z0eHaXUiTlmbPqFCqxXu3y7wsBREF2
RaI1pDguslbZddecObiKn2nk5NvnRWhS8WU0bpQMXFBeyrykekUVqDmMRfioWonnpjCNu4El3HjX
eljHVJWH9eOFdtRSgbSNhxP7PcSH3HnZO8mTX9dXBQvccUesfGIW1u/vSpNxFLpTXvl+xGTSGGFc
lGW2SnurxXJa9btgpLGQ3z591pioRl/XSPp9t/BzZTkJwkajP4+iGQAEe2h25hQDP+3oafl42z0w
4EXxDZulSGoymqzTEniiSiYKT7N4X8yqtDEAvt9Xowvi9lsdHa06YY3CXoj4HxKdnJDyge60EG/P
Pw4120MZ69p8++VEuqIQauRSjwMTjFIYexjIy1YjKP2J5bkyo9r6Kd4sXVsIglg0uFsMyAExZEMm
Z89uMOoKJsHr7Q2Np61QoTGnlpFHCEDEiEdRa9+o6+SU8Mnj2UqUcIXio6pBh+DiyN46T4wrE77k
s2xMWkWhVT3E6Mrw7FFTf7Di+oArZ80B/NLKtwGvUrc+5L94ghXiPCS2S2CkqbA1Z2wi/WZCbIYJ
JENCBUDmk+lPCd738jkgZ0RsscGLYLMs9QMWJyTkEkWj3iEgMu6/Gnf1Tk7uC536BYVK33GNHmFn
H/Pci9DcyrRZQ1ur8Cg1cIK6aY0gMyxRR5M9R8vmWaQ4+QJSOkGGt53FRd5qgcg///hN6FSN4AQG
edj6DaAsLEKWu6XqQBjOAtjPHyFex/5gWfg7SNVXUJW2ZoUmyRXwc0uuXsGppFayT1t1s/1mFgYK
ZleTWLwSD/Jza3GsS6Gp94nX8ed0HMuiqYSU30RiH7ySVcpbGEgxBZ2JKBIBoT1QiTR1xVMkO9Pf
F+ciLedhikGaG7/Fjv3XQYUkERiv3ifrDQ0U3TNDi4rL5LA2+AgbhVONIhlkB+UmV+n0pNW0vW1S
8Wke+6oU5OBjgO21rlK5oDl3ONquR+ux0qzoNNbn3tC+f/hgdVIwg9Uo8Oe4KDcNyjFOGlmxQN61
ejcZG5EacAaPa96MAqpI/uyfGXD9HFPx81wpDedwmaTn9HstTikPLLH+clCKC+wJ2VGVP1X04cwW
t8qa5toEIJmcugPbLLceGczDKdWa6jrKew5s7Mx3vpphe2Ok5KcHnwB1c3ouip9yaHf4o5myJS7N
MSJGTUd0zlCL/UqrlsDmCqAMRqmmdL2HfIRq3ibPuGyHzx5I0bedteImoZKAQxIfBQVs+oR6wSMU
8mR/9uiB2sGQLmGWqF4MpqRkFOEm5pLQvVVAoCf4P1rqLMgyiYCXzbqF+x2Oyw5azo8Hzb1xO8EQ
iRJp5SS7Ev3MhQYWRZPIdLzvZdWy8Z4qIMDoOqSqcVDAiV8resPIYEVEshkaOv7ChQdTmFWbmyvE
yXQ+JefpzgK6+GpmnPCZvx9hRiM4AnDEiKkCRK+g45qmOH96YNRm9eVEui4/8IYLoAlew9YnTgE0
CwF/UyRk1jYscAdrC2P2ypLgtMiKPAhZPeFpFAobj1XUyAzGLgo3+styZ/fVcl/q6efGwo8Qucyi
AquiYEvYOYGBPt91EvKngPCVrD5SVLfTaGOjmaVlyLD9zQTwQ2korB9rSPZD25remFcGNILAUgDs
PbdI3hQ/QdOCeNX0xmNG9CfZeBYGWbNI7lizvsBhEk+NaWYrUs6Mr+GSFjOqVRw7hM7wMTZwROe6
MZFY392bg60TmwJa/MKF59dfbIVlDN0AyCKE9g1hpi2U8ciiaTzawcD4h0nZTFrpf+MRnbXL9OIx
fmH5nTvk7lb2wVa+XcIdNq5I4Zt2KqKsJQTzrqqucm0M5UocE1671ukmWkQqy2Btqg/Qr76vxUYI
9VaVgOPmtPFm+LQ6l2WSg7DF1yja+1d5EIGT6KNs153Ow0BnxiCS9rx/WJ6DEq79lYE+eKbYA0+P
PnAJFd+xN3kcZdLKGXs32Wm82vRyHvl7AB1yvVjuI2PqmsoaI/ndw9tKpR2tcJXKeLOmcS+AmMw+
i/x8ukdLcLcjN1+wgPKieVIeNzQSoZ4U0t08yC4z1wTSJtpP+PPpaLjVBkVqxyksKeweTHAmQdn7
0wzyeQu2pQbtaQcnsxOqCfe9PWmiHE+p8gj0XvjQ/a2RjgR2JIpUTfT74FF5FLCKaM4bkHEcO2OY
6Ir63Q+1QCext3k0vgP2jNlaXDVOy12tzeOrBUuWlYYZmNx/W9pUasjEfB2H8FoVgWkRsluwHqJ+
vXwsdgrffs40UVjSmMGOhHCzoEtM72ozWDHC53mNhlBnXeRY3XVC82M1xwvaHxPr+i9QU5nx/8Jf
Z8kSMpIo6z/PM4GUXFrqBlZPKOqQWDUGEcXjv8ZBVULDfEM78aA+09W50EfwRRe4vHpGhD/OgZnm
K2UkiUEJS+/xh2Dbk3nA5wUNpe/GqBg9oP9orCut8jhsW86ELkB1C6VLArBSXQeZwdPmoXoFaoHF
Tyh6HKPFzEWrQXq2wSgQKem3TIxzVvy+pGQKyyNnrhi5WUZ8u/e67biRLrz2SXKdBp7SRuxh5Iyu
0rPMkJFf5SssMeQZNi06MZJPWj6LqT64OhhmhfO3vtjeXgjgdNCvCjT4QlbD7I4gBDB/a4Q9A6+t
k1X7v+6P4mRertMkBMKa9Pq2eJxNFe1DSR4OUShbeK74O/q/jEhM06BQ+VYylFwG6E0KNCdVQycf
LSm7r3ckp014rfNUym4J9lgAye9sG+U/b/xswHwLQfOGgaB99HbYRsQutiSJTQ7/eWulNg0Nxx1H
aDvogJdK53YnZIxexVzCR6YNq3OtJVRcjbpVzi/uIs3rY6ImzViiPiiCV0zWwQnXhqLXMr6RoRRC
rPIWrzzJ4olC+GKh84QHYrnie4kqIANFVDPeQerQPy6PDQm4BcL2U5ElpRL0iYWrihwimtFRXIgF
c4HeAKXtaadeYj7+AkDzeTn/Z7MnSa+hY7MP/M5tZj6koy0c5TZz8RFoglvHtOcRx+DrKKo+TQ0u
S8TA+fSVIXxI6Y9tWyF9DbyDsT7cNphczIUf4X0vhk2FxTQsb+qtcSQKrujrmHn16q6ZeJGlDFBm
bGg6NHWv/JKX/nPORv4hZ3nf82na8bXt3N/1EI5TjPySYJ2sIYGKFfySILGzjWXmDL5tmFmdKt0W
kElpbsbjU9/daVlK3UyWxnR6928WY+hR9DKz/e2HeXAM/Uv7v6X79/6CTAQV7cSBtZUYrUYFPQcr
4RldXRTQeWFsZk0eb+I8nXkXpIaW7yvztsdBscHWpLpmIuJ1q2738f2LgUsmfB1DWUejHHYhAfE+
4E+MoehRmrWYwXa7+viWhDzvDtj3q3f5AnFlDl7bwcuUY3vziPEO5sOQiCXwfm0P0YfxBN9cQ92J
jQyokE+KdkbDKA6TSkgcM1mtL3TI4xcV1LUMJDvevjIvT5FoAc8KkHCHCG2NMXBAel7kUricq7CT
ppzWLhAJNwDDmGKaMU6bazbgPeufp1cBdcEsWm0EOI3ZYg1ttGfzLj+laal+16vgzbONG9xZunWY
/6964BTrY51LpUB+4hxyzh86RzLI4BHH6mqY1QB2okHYg4CTbgLGJMWzjyyXtTlfV0W1n9Aob2Hs
KB243HhrilKPqrSY/m1caKVWpCdPldkYSjaQDM71y9UbYG+TClCDBUn6jKcwJQJd7LJRaiSWcKni
CsVDBfMEMzl0XPidN6g7wbwziKL5JfybbKNYYfdqWyoK4DOS6EIg+LZtrcYhZn2rL94hiosBJEPz
Ry+tzD3xCaY71YgT4rPvJ0xqlzbNtfP4vbEK/YKDXGLyiEZH9+17I+ZZWkrJjp9Wt91DM8xeiW+T
FLt+GQpD4joKy20CUfQ3KnIlwKn6eZoVf7o3VD8YsMdXj2M/76ORC2hmgl3kJS0Y/JdCqe4BIGXa
NVuoVvPluROqKKwxDR1Bth77b7ffVLJLdjlmwUQtJy2AsTi0t2flXQLHU/Sbv1gL9fb2Rnfpmg6V
qfRz5GBQXUPF3Nu3yFhhWsBVmDZ/j4v7B5kDduLdPcfKmmLCVG9qNwdR2219kH/kYzYDdCq85f4I
qjtMUPOiOW4YUkMR2QyGTvSvzvYHYNWDPcrO68o+Jsb9up9AK05a9PfEdV6KG4YCN3TATyhQSWUw
xYOE+jV9WfTbrKNbSHWQlTAPCWoV4OxYzatpQRWtmjmEFeAuwKWoTI3HKtJQm8IdJuUE8MsZZWjk
AxkxMMoBnT+aaCY3lNARJTZXnKExsAP7smFTQrDoknzbgvFY20TQn163L5c0HT8am22UMbRwWgMM
l+t8u1WGEEYb8fUm+tEKJSmoV6lit4tcZaKHMEmYVVX25TADouYOWKNgck//X1gOEONPPVY39Pbe
QrR+PwfMYMUKk8eOnz92q+DEz6aRVqcM1WANUuLzI2ab9TrGNtkvZmMy7XikyaCBxuKD6bQSFgkD
S8N1TrpIV2CUnWuVCQyon8/w891TK3rddqft0vPUV4AP9vZx4CqdNhlIu9BcffN+xLVi5TbK8lI5
r3kL380ggu4co9IUTxzWnECfJeFxBwCvOa5pvVsNXg/VjyfP40q3eMxMRBtXieBokKt+OR7V3WnU
A0NRONbdwclJ2ntTPUM9OXrXh4BdCd4ZoH8GoNfiAWgj2s7kOtW9un9EXv9fjTCroeOaJl/8X/hx
vPYyp9bs4gSmLm6m8BF7+TN7/7zV5Mw5MR62QVSHPX3pJVKnlE2iqfC03fTIyOwT5+loqARjd7Du
MSs7LXnwtpv7v7WDg/LNGSZzH+jsGahi7jrFrdwbVrGM2RT7bFmbJ5iMGTfiCMf1Qi5vlwPWS9jG
XbyjJBlRbamJaxFCe7a5c12MTvj9ebp4sSUTHy7BmZ/saDNmH0NUJ+jaG26nwwEnkTzxGyDv6aEB
9+rbZbqBmJyXLlriUzaudB0bhc9G0hzU4cPZQzq9WaNlOzIuc9c14z+SVmH9BzfqSshzOIfQWhdY
AxetktV9pYgEFUTrwfRfL0PjzooCniZVga+i6Vf2zgL6qjffMwI9PLpcvCjkRM7y65HgUVpgEVHI
Uyt6cT2ag9dY3jvQ+HnbY9e+Jwls7psWEWgf0lMok+Ykpc7ZVzNqiVSMG1GXYOk7TIrBL2LkBDBB
kvjDIrZ54rdsyvBFS4OHEnj797+OuLaw8oIwTr5naFj7wsWtRfsoFw/4ZehsF3OrCen0tOcOXCTl
lBTnbcjS6NT5zwagksTIVp0cFrRdriQUTYG+2JosEp43REiq85xmvhGzmc8L/7hQxUni13jnlOPe
elNZCF/BlF+vXeTetXU0RA+B6uFdlumNz0YzZhb+9M6vYAQm1I1kUf6f6YmTwwUhUYBDeTMjTXuX
gzAQaz0QkuxAOfb41YSjOIcUmipF7ByvmVAmrJpRvqSNbMbAGdiJ8Ml+dOA/abthV+Q16gFdwDGm
Gbc7ULQNUKYe0rwx1mEwVSaD9OV6oacvAjKRE5fG2Vz+HKLUU314o5BmDRIf9dCRb3z06pISj0jJ
UqNADfMDJ4OuKUGFROp6Xe/7sNK5HPjl7p32zp38s3GfJQ9VarbsnovOnJnFbrkznkWmhJYowkN/
IgtIi7bUhf+k5Km9NkpxwLfxeY6EqMwKZ65AuokC6wJ7wpUyf65uxfK+bl0hgBC0QPOvfzwCBPka
El8NI9c+Tfmmyg864cLJ7GNwwoMgpqybCJdYGQ7FVlI9Ern2gG7ZYOt5HP7d/M55cRK9PQ+ABfKi
abrgPegQ2QJqhHgdeBqnemfirMWsMKXAJdSXBQso1QehVwXlKQujTdFwbGHjgwuzUPNfeyUWh4Zj
sTSyxRrcR8VJ+HKvz68Xvjq6uIVYgTyZYOU0gJPr0exTDo2GvhLLRE8kG/TG4RXjMj2QF/oz1+Ze
T1BfHFEYCVd9h/A/0VOEoFwe1FZ0tFbMCLnrLPLJ6shEXyLOPH+dqfud8+wjyNHKeai6Ms1/uzAR
OJP1J4NRTgKonc//7SG8bRV8DQR6tmk2L+jRt57MnN4L0mFnXRv/SRGFMEfoSZe2w3SDj79AkuZ6
ovSQuTrDaB5zpxPiUIv09DpVMsNoh5dhbJeX9WU8bd14yYLaoi3JAr25Ui6gcmhZtsO6RX0bxjDE
7ByNL2Yq0Br+7dG/hSxhW0FbecvfeZyhwLFGonmVaEDBTC/iUABXivLA/tpMGvarR51adxkAxH2P
VTKMcnpsi4QjpI6mwDr2Sr40Dm5ArbWqACcfYP+OCxnQAsn3GSPbjQ7ynnRsRHHqBg6TpxYRWHvC
PTMriBZ3kLASlteeoybUEkzOe2lbO0bC4yU0xQZKusTnlIOb5rMx4aiYb365opFCs/PYSxtbvQCQ
lKlTuQd3OEmdmbV9DoFZX6CZZuJgQQM+jxfkSS5JgLQsbWAEhBmXrXSU0IC5PI9YDuFtxm8OaTQ3
Kmg3YLrqIuLbHqah9QGjxTS4eoxTVnQ+39wrrP+wwI+9n+iKVrQAdzKfGgWqRlDNZx1n2udytVIu
t6DTNVupylDjQVvlEvC2cr16Gq5QYaMqKAc/hMZOAV9laQJMyhkmA7OWwg0UOvRX1KTUNnsHFqoc
qzpgzQegRfWA6pLcCAS8EBGvGhrB5PhKJa4WoBHnamHWGn0CqqjtkCcz8HUs5DwBGClUSvP7EcZc
9cXXY1HRcS1aVXHxtXJDAK+oZwvd73kez+/84L8Q9m305yY8d6fKy1O0vleVwwihfwsXBXxxezcQ
kL0spMWtCVTsQFltdN/FkVQzpy6TBaDfCAd1OZmVZFRr1fzVFmKJQWG3r6Z9OE/A5zb7U7s2bMPZ
7RyTMstejUPjO2vRRQqGK4TDVQoJx9bnNjf41aFPBYKX/ABXE6ek7U+n6SROMKTHiOJDTLqqFVtv
RCuYKM4C0x441EsqVn6wP0dou4FTj6bOVz83hyFviRt4UOblRzSvxFSdYvlothSqoS8xguyKwJKs
sMq/Ej7LKfEN/Z9QVrFaYYEP+36EPeuOKB1LVvv3XZWjVQk19Qf3tVuhvGt8CJBegktmmeZnpLMy
Y+kJQBdeqfV1Wl4Rg28EboLMQjOT636DamZJMek05tqMAt5IF9SxD3dAcfv2/0DiP3EUGI0Luutg
yMF5BUm/ll3Y/YFRb4TfL0uL6s1nASiXb6i99z5TZwxxVGauvG1RgFS/TRvt3rvDDiqEzMOW88nJ
cwn2HkWIcZfLtzFJgz1aFXBAVQJSBoeQZ/FZb4SxfxTNqIy4KHbA8MH/vmCxsO3jGoqewooeU+Rx
XC9OFlPkKJnRGRxrD5UOympgx3qpPlOCMLBILKjZokEFsSTBNm+vz4p0SX5s1cNS2UurlxClvqAC
jMgvJ4EwDqc6c5hsWEWicqj1R/1J42rPhfanMNovAonOCZyfeQb3D43A2sHmm0SWVC/ob39vX0zF
amwZw7o0cH9kz02vC+obTXDNTX7ERejvnoSoiHrgGJXQqCGJNszNrvmGDuKDdTakAUV1F5lmfTVR
Wgj9oon171a8/4DuKyqBSa3k6YjqEG8FcN1gPl5ddMuAkP1z1j5Bvi66PXkm40q1YzbJB39pTvNj
cuVnC2vKa56NSWp2GfkKwTxCRLqMzaw8ejDnyA6KGEMZWNewtPEBX1FWibxidFtSV29BfG/YkL+M
DuobMNDKJ7VROiVY6Udu79Af3bHCW4lqBbS/AFegGz6sBNkU3klEJAnRdpk5hwv/2mebYmaavdS5
RTz8Sdnf20YcR5Bxq6w18QH/DuHLNnJR2qsRD7rNkNAl32xrN2n1CtyJmEGRytytVNuLXW9X6b5Q
s+EAMHbfbGfzHHETcAfiNjp1fpg0QCYcOEh823KCXWElXd9QeRx11GAG5SrK4p3O52dz1K8NxI+x
WuGAt+4QXKJkkizgJURcnDGdPy/kBQKGT+DincG10lL1C7Az+MAXcCdt5Wsh5BDvrLV12erCBmss
P4CIG5Tna9IydrsmfAe9dh0yaH/Fr9EwWDaCAR32ZTM5jV+D2aSHotaJXgLP837GhHZ0FvJu06Tx
+nLr1HDto8gCJ9jt0JC+kwGuFAnfUKINf4wl5eFRPzYPczD6qw+2bsqoezWWUlOqR0mxGo7OhnbQ
alOuOjje8TsOe7Me1vDGywqpb58F6C1NnslN19fxC3scjpF8/8VMv09PtPFiLV7e7iLtbC6OOCxf
T/vQQfZDlQ5jwqanqW2I4Ia3fPXANlAK0ZYj2Ip0dp87M8dmjqJSCYGlHrYCgp6oEnUlhqvBaCwN
qOzeL5A1fEBoyvbbQe1JdoHGNC2O5Xwb2OcElafrbGNCv/gUyvOz+FfKGfVw/oYhrTakjrGTmN+i
+RnZ/33YPGDNQAKo+9ikJbneDqVNn2SfJCeI40hDdOS/nTdX3qAIG3FulthaiIl+rbLYF/zn0xF6
oKJG0XjZMa4sUeOCIwmvrceFmWiOW2dS7Zm2L3G7muZo0U6BAw1az9M94bkBPwjudIGZf6S6+mqs
92e7gBEua91aufOPncoaKI+ubZJAZLC+afaVA++jy+A/hdHo/dGlpi+gEvH/kDVBBBQwqllxeI41
7Rkdna+8XOeZ3WEr69FwftoJl/jqgq6wS3u9smMSH9q4kKnxwVGLeV5CZJ4RWbzxrqKtcV4DwK1p
FD0PMnJXNwVh6UU8S+PDfQKucl3elBX7cYLRB9kXH2/5A1R9dP1ugmhzk0SoCvvoKLHajdHsikFN
7MI9GKbIs1YCEn+vI+h2TtcxiR9SYD1jRrrkm7vPAtKF6Yk/1yfrq5SL6ER8z+8Rna0OysjrCiQt
3Nckwt/rzD9GcEd+zDVvoKbVEej5EbqH+QaI31F9AOsw8ECxdWV86RsCGOScDgWJX5s1PoFYcFXg
JFabPR8I/lePuJlwgOUVk7+9x7j27fkZnwYYEg+t+zjoFpnNNly9/nFwqG1IrOhAgLFA4drgkEn+
YPMYP57p6zRLcqxO27zL2w2/0kRWD97m2wpLfTIJuNX1QT5Ujq396Obeg0rHAhjIfHMsxxQavqqb
lr3Y6yKNrofJgwpcZN4AwLyI1B1bwr9ZpxmIUzYl7amDj1HTsVV3r33m1fsuUDp0iOsWZ+fefuJH
dNNKfaisrzcqaIxiv7kOWTnqFonpZwye3y6ZzcJSMn6O6gJfoM8pH+MIYhJ6T2av2s0LNg+qe0DL
0YsGhRcxyzf8WfF13KeP+0Sl2TzngJhf43FUPjR03MVJRe9Hd48YJDTnOHjj32JwR7rXj6XvrZQb
G9F4dbEpOY8TZcDb4CcsZNCzOXkr4a1fJvm32nVzg0sf4K2TJKyYLM73Zcu2pSEwhOrOJNhg8zzK
lrAwmFjH2cUF0N5rKe8u5ExP/30ma6y2FAn4uEphiCTSQl3xSY+sRZZMUjvW5WkITFFxdjtl50U5
PWQv2eaJsovtG9iWzry84j9dWI2JCLOlmd1Ft2JQutYUjtIvSNqBhdd7TTJUkdLQ9HgzWUCEM/va
JUuSmbwltMKZWVRIvQvRiSsCABwqA4kvsoMbAK9Ybe/hYVHNlev906+h1lVwtpZ0OuOA0ZxkFRL+
G1z9qPqubrH/BQTQu8pC5QSe7KZ8ISjmQ1TB7jPOf49w25Jk2vfg6CU29N+N3QBgM85wl8w+Vwg+
JIJRJXEn0Mc5dA7I59uHDe1ANsNfKraTWIfWDkUi/eITh0awhMEAfVIpNV8P4UpC1I95X/kZEaDp
QLOQuutzZx4WvxORVcTRmlO+BYKUKGDN5rmFP0K4DgUcFfI3cVrgrYSn4Gf6XGJgH7KhgOugoEMU
jpjM3RqOleTdBtCXsn+tdHzwqxDfZ5tQSyJY4Y9isDq7h5wrLTDndrfk9MU9lbW6RVEpP+GG2lSZ
3mZkDeWLvme09uytD5oxq4lvnzZlLO9Fwir+sFsvctTW7R7BxjCbKfq/IXX0PuRwTH6blMiuTCOI
kC5PHQxXQJwb/g1eMgFBXwaaJ1enH6sj05hAzGI7Xt8UCyiZ5ihKqWxzd6SciwveZ3iGFAfCvFob
Y4z7dTbviLnbRaOs4DllveE5VjKI1H2Esan/Ws2crWHdFzezSFgLP2VZrM+QSLGxfuwxomWPoYU+
dACmvccK8esXDxS/qjD9z7tibTLSJ8EXsvjSrdeyWy/K05CQ/ybfbUej8+c3nhri/vPGVDbjPe2A
5r752SSayLpZYFXCDR8FBu9Id32Bxat8tHziruzeukqpzgpllTtNlmaq4MMqZN/F0dVHntK6o/cA
9AvHYkP9JeAXL9KvyjdR2T6iIs7nnqSkzTayRbFlMQXB3dmgxsEf2AMIpSwUt+x6di1zHuJNWwep
GjKaIvzqTrkBjR26rq6hUi2RMKf2ZHX4suh/bv+DgyMoLJdVC6Rb+d07BpUekYmZ2xWQ9JQnxYiU
LqzMsIbuDf8SGjgaigP6Xzme5eh/udsQ6q2gwGTzBpIMW2ypBjNF6LHHmW2VPwljuEoe+aTiYgTd
Lc7hJFp0ZYhRkvh/tiOFYW/OZ9nRhhBHmasxnhJoEfmrYvkKddEBS8FAiVDzRHWFDWzkc4Heg7PU
ZEcQeOdb3MSHxvwNUyO16tuk1VlldmN3r7MvgyyiIPUYC4qMzbOJRGc2nhHCU53CBoCKj1Avx5m+
qNG9+lXOxEwfdMWdu1mga5Hh8VVQbHlwrHPnulLOTQlIE0Ui9SfmmLlhw/X+oDICb0cS3TKgiVGM
t/NjuxyYlHcbO7iQQKV6brQFTbcsZY/JdEFUAvJXSGRFf1i8aonIrDiNuxFtMSuEaL+4XpYRBxk0
Es061SgdP+DS5Lt0BKm9Vu6EX32dXk9Arj4aPme7nGl47ZPtCpWvNEfFe1NmsfYUPopD8I5Dt8qY
WzUg9O5pZpAM3iuwzwrcmpcbFKBvbP6N1TmHCG1238YOAmjzItl3+SrRW2bWC4ya4BKsGaXUyCxR
1XAf6uJR1WUHtDUp+YJSOON7dWPxVkgwirczlD5H5Pbk8qMXVFOIOww+UY5Wy/y0SCbdpKyWdhtG
fCiAVtkE3ZCf3+550weLFSKP0hEEIzDD0j69NCIwdnsPupmh0GxBRTcx4JaB3ZDXqXWJKCJTrImj
TDheONbY2iMMhAapWb7uCQRt0T6ENhwml1alxmpZSlnUIULpzvBDzRZClClcU2H4ZoEXQHsbJHMc
z+tlLuIUJuuL5Z3Yc9Not+beTloqQV3CXhrJOhLeiHDKrDeGSlRIts6y5ubxltbV+TNlEfIELQeY
3p6PGbd7wzYB92Ulc/wYsyivLgtkVEukHlr7mx00LH016cjgUDzGFJYddWZdmzXgd+/1MVLLvoun
xyELNsk0bnv0ue6MKVw+Ndt9GCccyWwVqG095OJ8sppUgj7Mg7GU6701wSQasVXcVwFRXc3//zm2
jnkq0RxxWURg8uNsRomxUHDjyr15JQsUEp+hFuhmTz++tLaI8lppWDAWLkjsILPi4bnhus3222cz
XBe2Auq0NsQEFeuL3Q3DO3Y1py4925VgiHdcm6xaJEpoCOMsKL/qwpnGlJ4mVp0IBOF6u/s3EqLS
fMPM6PvQBfM8gAdcvxKbHuPmBlJ678oLhViYKxmZKdWInLceKhnvgpVQHjYeYYSO/w8sZBZeS5Eu
mDEdTyDh6T0dYWfNW1/tFcjSuOcSoNSbbfJOLSLSC5EnWgRvrV9mzxIHKwW6Wj9yvtwabRw11msr
zmw399kTXzqk9cIhcJpuB78vW0ipJNXtR+y8xpETwau7SAVq3T8D+djOj4KbbORLXBPh7sMn6YGf
k5u2z0uNdIxfLIRBJ8OlfBWy+67swrTk685kCuV8KVk1WoooRbidQ7e55mBXokAexA5j42ukWmic
Syl5ylhLg7PKSkuUAskaFN2p16SIUiYVhE2RWEFYgN+xqD41zyVsSK8w9+F8dgI3QqrFExbREQm2
IUkSjLxwyzf8ITHe2hLw/9t9/Fm0e1Mkd8G+tg+AL1sYxQsZhFsTpQx7QjZZdLr9LOqQ6A1hGFkh
5NVS0P60KtGTF/frrLGeco5nYgCbEA2kwBDIoP3zc3rHQdfhsJDZY80FHswvEy5UV9WkjSPySlIn
3e4YvFArAHPgZphigrQv2m5Q4QDKRGdzsA6WQt+D9OJdT4Xv08g527Ux7aPFY9kPPbk3+3Tbm2wO
9RnY1E4f2p/ixLj9JyLofse+s7YHG3X35GlTDVgnBlMAxE8iWEE54i++j1lDd9+dVb+fZhE/bNNU
/ffdClhxsjQsx3BTxd62YK+151Zy3Kfg5vikXQN6yCFhm6JUjAvHI05WiOasmB+zVV51aFnBqyrY
q4N3dzg2cVNdSrGdmAvrZqJ1jVb8lkdRJ8N2TPVFJdf+o/RdNOK88VUVpIch/PGR16lo6iAFJLwL
ExJmCiqg0K92KOZlHcy7Mtd757X37RGiyjB5rqTVf/Bod/XdGYxKZDLRCFMw6ubIa5upaezCHAEr
I4x8j89NOItMEFn4X2ypjVSwJhaMZOW+P7GAVIdzA8hWd6fd2Onu4k5EeQZ8FDOYhIc6zmKAEGdz
EF5oZb6gc8MTToas9kO5SZefDGQgKjsYicKs51sjE19OgOxQISaKazwXPTaIW6s/fB0hX1wYw7QZ
8l9PGTOR8fidHl4jYYTXrTl+j9A96yoVnbt8au5O3QLl5jQoAfe5h+HA7yHC1AI80PSBxkAY1XpO
a8oArNTasQjTYl4NjnfOJ60xQZHbig8VcCwMSH5XBD8EfV1hYfzBLuJFSZzMpJT80tZaq03KOBGq
UXbEb+/d1WEciHgT4a1AY8gU5gy5UdKl2Jw8iWEtD5hoW9kuZngvutWefMSj+0nZkjIu2spiot0o
siNj2lFcyBAcJZPFsdSD0kOwdydOHYhky2oGfvYgDA4+V4HrD48g6cOdLn+dDoUp/Cr9xYt74Nat
RRvK7wHin8uNaovrTmgfW6wVq1I6bRZki1KUhcznSfIBV12LN6OhazdvLI/8Ook/iwApTVpA/xfZ
9dV9uWBw5HgnR2R4KnQkj8Zym6d1PWCzMMufQxMjYsYkvgkvNktiJCBZTAdrce8Si6wpz6D8kFZN
afLloVRfB8DpWKVBwbxo2gFwkzM8/G5kuExhKrnyMAX3E9J34q+1Ncq43q3Y376OB0mDfI/AtasR
Q93Id0xsFYMihLqvmaNpbZfkG6GxeKwusImkyU2+i3bbdCKbfySVqORKMywVivEiquKfUN5AN6e4
G2caUXNQDtSu/NXD67xgqIsSq3fdLiM7Aw/bOJomkMOr0r3iAZtwXs79qbK4W+JBEvTsYgIIPWL6
2mLi2mZHg7PVM6VHvPderNKxTXh7evidLkELh+JFY1CXg5Pkl+WS+b7N7b+toe2+G7h+ZKBpGq/p
JP5trCNmJ9ni0kxhJbrAG820y6XOSrzfBojIQOdIvEG0A0hto/Hi0KGZsV2U7erQKbEnnp3bTUyN
z15AJ44ZT5tGDMOux3vlruKfkBwaSiTCpb4j707b/yBBw2Pa+TQel55cffjdJ17UylOS/Ub6349M
jKfa+HB4NYj9ppJMxAHsYbpH0j+XyJuMZYOlfNOtWCHTXS3nOpQqUjDO1/YO0FnaVuwWl8TbeUYE
urUs6l+W5CTLMUkMeutpZpC6snomwaduYCYv8Krnse+ACEJf6f7E7KMqyTycyKhC9qxFkTeLB0gP
u8Ypvf8jKi1FuEwT11lBIcxZk8pBG+Bpax317M2SC01TaD86IKUxwxtP3CckaURNFv34lU4EBIRk
t4Ut19iM7g5z/2c8IXt031YPTO+AYX80hepyhAvI9d6zxoLPTBVzy1xeNkNeyzmsZcu0kRQq84AD
WyxczqgXwLumb+kEySfvDFPi802NK3Ihtq6uDbX/qV3wwTTj9GMl8A5uJDChJAgowkKpwoj1cGWF
DOIL/qwDVlVL9ywWl8RZU71It0rdK19CpwBXsoXVc8IrcChrWq4OdoySOPdTvvfWk5gEa7LwcSCp
v0NVq39ch9HQuYdvShMxvMUULo9y3wri73SXK/hu4FEWRu9jnTrtPNoY8NWQjhl36pz6I5RJC+Z6
qMjor/npNSlFsdIFgp2OfZChjXXUAjF+phUk9AH+KgpLd4OLxSEDVqptLdhhRSNDgkAmrcJuJvo1
HKJzeOYYjsRZ7PkuIi1ahOtAv4QgpM7jAnbSgGMPxPDn8xvdSWiM4Ibof23NgG7wd3HhzEcAK7vf
GqEbU8hfnbQCUH2DJE1qWmTowfkJmns0bL8s3ZoSQcyMfDylSKtYBO/K53YIDP1vM+Jf/ZQUiBXP
M7YviqpvhTbKkGqLdfMt+jAQK+7hLSoW9/Tc8Fde7TUP19XxKrwo+xgAiholCWxWPeFNoZuruDkB
YX1AlWpUylF4ajU69LWZGO6BWwMfoTrs1YFr/4HnPjMZdlT2XWeki6zLJCzbPJdKQny8idGg1Sh1
vdImn70o04eNpNKQDO1beAKQwEWpu1f4ygPi+Jgl5F9t3CG6DOEaC5+xraPsiY+Lc1uqDH/HOqUM
gqMM2INKqwMBEjjLnauyVY2AIzLqPCdPCngtRx4s9DxpAIiO+CTF0pXaWIcFpoRTIeWvWPgqkGy/
S8HTDdhGIqJR5ToYXeRNfbOdTDmn8vo/Jel1ZmE05mp9ySYJyUrNxIrwumCTdl2c3Q63ORy/PTtV
iXFnk62B6vNy7UKFa8VzcGUkw363pivRT0y4MOIETYSLuCw7MsZ0Cfd3X7T0Hhz2+ASnTb1VJt+t
F1rh0JhiRCPtJ6SN7v0uIiNr7whK5/dBPc8WIy7ze7ziz1S9vKv/yq76nf5k5/Pv6NHfk/1D59gM
Xndm0NzEPjPav2/OLfJMRos6qspCRTE3jisJfa4R4a6c+eRB7addF/dFNhoWm4YGu71jt5ywlel2
ZQxCPT19EcEiAtEpjZM8Oa37tLIBJ6KaPpdzTxl992npeKThFAkpvGEV35mVV7XaPtMQmyeWwBsj
jAiEu2EP61DuMCuCGTYVH6xwy6z9eaDOwrwpSErzCd74iImfQkaLrq29Nw0nJFQyPOdMBdREHDE+
zpiWkxBb6RaqFsEdDyTrrUqE2qXbZCJTVoCsnvwfrCuda+RN8oTV8kJ1zGIkkZ/obHmGuPua/KkD
ffEtlYBlfLmc33q3CBXEZqkPd9B2lJU8/lr3rILF6w3cTqpnU5mYrjKZ4qw3ivzY9Tzs2A0x5uq8
wSiaFpF51a1HxYVs8F+CHB9BBtCjmMx+i2X0V1aDNZmXZ+UuZUQj219gANTzTvZ2rW10wKO0o6y+
CY9PcOFhRVHM1Cx67MqllrOxhLgdmGbUPS3NBDsJQRhHa4NH6C+INThGVCF8cKBkPSpyPKTrKzsL
mu/DRy5DaFRs2RiCOq8+RkkdbrwBM+Ey+QJ/Z6dZRFqcinlMvGIr8/6SrBvuECNxfKv1jSU7pId/
SZA/yUfkwBbg2bR9gUEJ37ofbbx4xFwA7QW/gVDXAEbpRZZQGjYe4u61SwF9rN/nXxXFBxX1hPH9
iMsjb5oSpJdQ35xwDtFiIjew5RUbv0uaA4ubBewBuWSMRWHipSK1X4o01gL38afIfCfXk1SM557b
PGTrkHR7b9dQ9TlLiygthtDqrBfum14SePuWsV0h6sK1qqHJmphr9Iw6kidWRdcVrzEKibsTQuun
31DiYDxQDSaSVbr91ZCaRSusEhwZiuVZ8M+/uOwLCRmXK890L2QC+BCR22yUSJ6+jkIpU3jXb9Di
g7nWfawCvEBtP8/9J8hiL0paHpJhYHEvbD+32RXzUNcAMTX8z+tYK8xzAPwuwMeBVJliAytGWHwl
WheK6CISSeYo9OEsRCJmqmRVXVwbk/l0Uqh0oHuzRTxpLxdtVXYtcRqaVeIHAQTrsojjfAQgoyo4
yRV7UR8QTvMmAR+g4j1YOmqR5HFw/zGzAiVBZoXEdTG2ukG91w0LMmT1yA2DS6ydGPtiuYksJHiv
NMlD+T9pZ1qE/3xMEpSelm33C0hMPa6Bzp6UbpezSAJGZauEC/0nrsNVfnfqKHCcslrv7VQ9q7do
iIkl1LCFKz+bY8ulzFD8hz4gfIswToS+p3/oN4vXaBC6CcnrPhxfTz5hBd+aRYFVlLUuLIq3+TuI
R6YAXsk3lHjJwUX2ojTQLrn21I2GJ5R4XgcoLl6ZiUCquIsln6w1qoZHBfsDRT2wGzbJeeMJnFnH
78N5TlZQHXcTCf5cZ9ek0PiNBXYT5/FHRo6L8iwkMhBxMte/l5duGbW9kPOWX46r2O3cajjbMjej
0gGhzKS+uj99I4vflJhC1U3z5zEx/dvV7TiEOGuadUx+JlkFA3vi8ID3q26Z3Dz//3n2ZfZ1TFKd
dAexUwnTR4C3Zp97iQbjq5hk3czNvH5GoPvFO5mxUwCODeTZ+pDBq/LW5esCpCTxwP/px+J9BkES
roGDcs2Tv7RA+oiBE3xk9BzNgJi9xksGRosuBVZ/jcgdG4lTKenmCO3gkWyC4BxEwUrkkVt6LrZ3
MDMU2FhZ1rFy8iNj54/1NGCcKRgKjrfRzLK1K4/ZnbwSCQmLQ7qZoZTaiXOWRhfZzIA5eUW+xszs
UBA5GKJyvQzMbEyzPKjxTh10vr14d3xH0N+Xh7vAejnJSb0a3QKJCe6oxjSH9MrV/Hs4Ac2rHgGx
eCp5lwJmd5PdHPEpn17Iw/IkB+kA6sfKeSh7GalwGTvoV8gRqinMCLo4RI7YySezA2QHBMoYVIM3
/O5sKux77JUbEXOVmVCZoyinjlsn8A+dA2Hk0a103stPk/6pDMuAEfPNxTfHQ6h2iaVZ3LsggM0M
+NR046ekZy+FfYF+WPEqfzEU2XsNUzG+yUJBa+NIuIAVO9UnC9uKxEXptEh4VpHQwrCTpj3q7040
1khMSdTlLvvsC7THWEDnaCFhIrZkjcOFI/rqEOfgnxPa1P64/pPMoFbkdOj13/Y7JutuJedd1kkp
FR4z6ptsWnAkOLm3eb/KGiuBd/71lgIQHD0AXFx6hsnpruRXRSAgNYIWBM4vlZkKMnenpMLao97M
7Lc6w6yGu2bMSHdYl65jsDQy9lKIqNwdGaJPFW492SoUFW1WXIc8lnvFFD5NE7X0FfOvQfS965ks
FbpYcEeumEhqwhQrP+VLBHPQpBXjG5k+EESA24fazxl7w4YJXfE01raW37PUjhxJmz+U90dXPbYl
YI2itkQ0PmUj5Q3z/JFwJSgeCC5fK/uz8Wyw7+0QNzrBbrzieJbJi48/GEiK6ORxYV0egMtQGbYD
GxFM8c+rwq3Q3IIxq1DpW4LquxDSYGnDBgmWabemuKklMN6HXzOYv4AVX8VCUb09TK/QF/t5qq9y
7u90PoW72NWAZEgb1dW2eFIZqLSFRk9qIVdyBYsnhcRtqMX8lzoscywzFcTmD3qF9As9rWwX4PKc
pF7yO23YbYvU091MeccGbk48AyTRfWxBoDZ5qSeE8BAFcrRvhmt0J86Zge5NqhfkrzTqNX+RDOjq
Mp3uXP3afa7z6wUreKMc90nRlRiIOOe93i3HQ8HXW4j/DIbTccaO5j0SpC7mHMEnjUSg8IF7PpEw
nopiIIip7YQkB5pDF3S9ECLlajx7GZNVsnSPmLJVojlbN1rq0TGYSBIzFmFoITt4xgBR8nEKwaRi
M3vcu91RZR3GyJ3swjWYHKLxteWCUGORGVxzqnPqqvIvIES2UCesnbbe0trn4iNScxdTEJEy6H9/
qNfanMC6vlwRTIotDNhXiYU2w7m2a4wjlvukXz1hVPWyVEUTB9thIo0A2gBFS5WsGrqDcgj+tB3G
b7XwMvf6Qnmc0P6CBS3U6nhtg+jUrY1Tbkjs48dO6IakupE4WsvcFadDw3YiPXK2ZwX/EMyDFMGN
Ed18TYegz2i6rz2rCgE8BdzDv+NSXH+gyKChphNTg3qn3BOtNC441wyo6QdXoKkph3h7FPcT2p5w
JW7kqrffhzJwqW2M0czhTwyiCdFDJ7mr1zpgSiHYjWECyTP73chJYJd89TbkpndBrlDjrFIZIGMt
ptwX7ZqzSwYN9EIgl9mIU/Vg2WtzbB1msBsH/5IdLkJw3xLqEdGqJDsYZjZmQfeY7cJTXylCwOUb
QmhUxwf5Dqugqwc2CL8OGChoDW/IVwLLKKN0/q6Bz5W/jDBgwH+1DapsYhId8BrBSN+oQDR0OOU1
aPz2BkE5RxsD3cZmvqDU2/kbWf/KmSJEUpQazQQgsRiyDy+V7/ZGpmpKux8lVpeRE/bRJ4rXFCCJ
gvQFvCXqTsJfVfAEGrLjxA6Ey5V6c1eo7hFBs2WRriLkU2dB4c+GtRIYIs+YjNqaCvlReCY61VYJ
QElVu0RnQ1/wLqdUm532R2NZp8r13VAuFJS5hmGfkkG1F2DkpvUjxLWfA6iJU6mSmVCfGQTssOPb
hVAxWfxbs/UlhW3q2m87mS1YIXiVb1y+178fuxQ8ferLLn5Nhqpt4nrRgpfgMoD6tL6MaNCyKHRH
BVtEIIktDMQ2NtCN0Tvrt8ZR4wqdGu+IKqYM1E/aiCgjv7vqFgqKmXUjs/NqkrI+kaCp3DhG/dIT
CiPGTDtgJ+rL/223+g+WmTFnL/t+/m28vmlhAgk9Lx7YVctn4zSpCr3HNcRJrWRN1tdlcGHKYmdJ
m7MNVXY3+jQ2YPlZOAp3P+wkHitiNe/IpspqqBX7wGmEPoThiIp2lO54AboCtsSTTKgx0GKknziI
kqN+6IIEvl7cmWjyx1O9HpAQ+phnahb082FAb/b+32wgiakCQATdxm2b+mOAzwbLG//kLpSQJ0D7
HbgYVW2QOdNgPs1LhTn+9Ks/fyg5P5xAid5j9UfjqlwZ/I4ulirebCwB36FKI+E5r9H1PcO6pkp1
CdLZhSWaTPPQwbquE9sGxpurPaQezEREyVQbYzeyvq4eadLxhxxqXwWKcfYb7nZiDbex4NoY2iz4
UUWtN51dE15PA3xiQHRSzCkLgt91RCNMCLIkb0AvSuDvuv/49NIvaygnoNdcZ7bJZk6b7biKmvMb
UHy0SdpZaxAx3kPbAP1PtCO4EdDcutoSSQKA1IWgg1QsWQilt61robNqNQbcOzvGF8XQ13F7KXIk
KkYcU56LnKLckhu+zWsMlfbTn2ckogOoO4CLaAMT05wnui9jv1YauHNKMZyj5vjrQrKjIgvhIEPq
D1uXDZwCyl0D0mR5Jz+RP/xFkJ9rOBPaYUJTneOA1fF4jm5M5OykAzY2mpcXNUi/NaCyPjDqig7Q
PoxoO84Cuff7Ro/MmtnCMK5Tct4BesSAoyfH4DHDogrWw99OnTmtvsAnd1whFY7Bf2UvQjs4L84M
O7ocApGJcsN7ylBZm8bHLsTobch+Uu5ylOAfS+x+54zk+J95zKu137aStESL4PqTRACRygSgZDEa
Xhe/h5KukFPNdZ4v8XFsRzKIFC+H6W5dHTtpdGt88JrJy5j8beGrhXD8hRgU7mxq6DoRhfuq/pn2
mfwb53lvI26Vltnkc00rvt0OnnIKg+DnCR6nmCUZc5h3Ytc0bP4CNIcoRmDoRnwL6oeb+7dtNIln
4C5YPEdsKkge7iJidzoSARVzRwGv+MuKBs1V4VGPyURxk2/fUbx9JWILtG02JG6o2ppD7nRtVjAb
drCuGqBLoiba3I2aFPD0VjotMUsYSVv6i+GtczL61glGyXupKwk2cqJBRKTW5NmO1KOJ11uMs/ht
TtB7skuDpLeFdvSW0tNRw2dvomN6zPwa4mNsSHh+n1dLe2YTFlSjWDQCuL6NNyiqbpjPyZeSexmX
2r7KIheCoWC2EbYQ8SiHo8FmqTizZ2+zHYRpjelGoLePxxFURljLYvrd00Yn6eyDVufpDgCcsI0g
7EQltQZmYqfOePx3Rnjy1FypsEF7wXzME8j9577CC73W3ccdRgVx38NsRCSJ9DcWkkCv6Suv1h2g
rcsaAe2qr6OQ86jTBGGxCOcnW48+eApFZLLyqFDaT416wSxQMPNqF86tiYdaiw8527dJA0bVo1pl
lFJuGm5rKN4qWXdCP2sh0drZgsdrDi8ciNxBcTWzTEUCbwAnoaVsyFuApKxX2YoPiiJwpZA9GBBt
f1kSnzQAadKeAehK5GlT3sIl9T58+H3MYpwNS1th/scKqfO/05LB7EtwaI01EnEH0WnujsDY1B6f
aEtVeIb9KoxZOp9XAigdaTKJKMDInK1cYmWuJQD2ebt0LhOANGnzVDpUCvJB9tUtEDxAV5uuzPrb
6WbPWZX4eL5nZfYT5c/o4G50h94Ab5E5HynimYn0R0lyFpJiqJAcqtHJrwJYDUnWAXVyw0oQPOs+
KdmccHjkw2ur6rd+lPyl3LmyR8t8VGmuaw8LHwu5MgYbq2r2p63Ccr9kQ6IO1ne1fPiEkt1XsNDT
ltoWYIu+vPjDWgWR5tUtTPNi7SqAuxzo+L12niEkhSVQDfCwCNG9LSmI2LZf8uVJGFyjdaYrslgS
P5MRTbMPZyXjoP1zj6hB/HbxbRRfaQAx1/+8IO+putJpD5YvXcIN0kD2oieVrrKpMPPO9iAIwcE6
NFeRIYSjpk9ratoFNhl8l4C2ljklfPl9cQEeun8++W6Ju+trcKS8oSBaUQ+qc6qtD10k4yt0JfzI
vyAc86F1A9/TOsbamUZ6osn8WE4v2UMFRlyKZxcrLPJ73vLKV8QNWNuHHrekijYr47In9ggxe/iG
yh16g05AbwPKhEMT/j5OxJW/3jHbIBukH277pgI5cMcLOvFOLK1AVgLT0FDQz+ti70+zIAeN5l9B
obcm0jmPY4S1F1xXroMbP3FcWX0CefKvn/dC8tgpMOkBDG2UvN57A5kKj2cgIWz/DXdhLWgdeXAw
MB6lPo+tLBwe5tKbaSof+9IaB8Qm1TPbP4WSPbZdrF/CVfS+rLiKfMwPDAgxsgWQT/NaJZwzrHy6
KGGHIoeu4Q8SIf/SW6eAYIKKJZh1Seb1ozRIH2dpz3NA6ToUORLGyiymLqeNdAxh8Q/zwa8StcdY
ZgEqaHLxp/BF3xu37LmUUiXdUMZj7KaT08UpS71oWxEbuFVFY3AgD3pEseo8cOIo+oF2n44Rmte1
OL9hQIg+X98eOWPlhg20sjTcmMedYLcqoTjhc9r8K8gHad5ZvO5N6ypCdqFBpfl/bpIICUnZTKR+
w1IrdyFHeI9togg6tZqVkxlF8mG0lX4a7BI7z+g5X0CpdGtIfzKmL3GHFOTxYxmgCEeSfKacHPhM
OQIQsDPMGaf/dReQbSGr8Pvg/jILeIc4Caxd9wU30W5mC7QcAM+MjcHKoy0ivd7RToSsuHsWGlbs
1LBVRbW2EAHbGEE5dpqSiP6vrfpIvpWBGWTTzKjjtZMq0Vsc/A1YECVxSHYxWE3WACmZrjDPm55H
Rsl17B5oAvMcwdEx36Sxz4ERYOTchzd5aoX9o9QvrbA63PsuBUZLh7ttfaKTLLxlCR7eBo5ehgY8
A0TBT0hLYNFWu6rnJon6JbGrp6xfhxG5S1Zec+bmVUauGb8uagfOPyasYhqbD/Qqnp8Ipus4f6EP
oMociVqRLl6wX2QpAV/iH+S6JOWZYg3xOBKTZUxq6q0oaD3ES3AZcu+JaKLgrBlYzV08hYyqNRG/
GLo5p69wAupv8kcBCMgKuw77nc0g1h7F9l2F+l0mtMoETI52IAaX1XZ+J9wh0RJ+t0rSosEKWRlO
smW2IeM2p4TOYWCWZjSRNbJpPiVVmAWOj5KvMtKZk8C1N5S9l6q79uScejFblSOC2WSiuJIq+on+
gOJe7Twt0B6VKubOt8LzJwQc2GU7/fAG07OBaanCiGvRqQY6y7+1r7T0QY5HmXtQKvFnFuRyR35H
c8Qi+O64p2bF0Yak+LNnrxikRQScH+xKiREjt9dmM9dV0dSg59HXKIbPtZvgFqs4dM0tiGJl7W0L
+LQAjgXQqw3zyRLRxMe8mbIUUqwjcdpNKuVTMkNy2hibSulAdTGkochuoHoPJUtjXP590QmTumhk
5FUbV5kCETNka0FV4fYVmoLzGlYewEgQ87I3WbpK7Pz2bgzWnsWvFcwJAPW2iZEzBUE2lPzbQywv
q/IyMEfRC/I4mdEGbMmrqr34p2CEoCilh+3ggHvOwXN9vxDjGfUZO/nxIIw24xZPKIZrjzM/CWco
lg7KN/HVR4bTOkS/geVLsQEwR587PvvPGQZJV0abNsT+NTepwCWzX2V9GK7XygjcwTTEoYg26mNJ
tEKv+SuZx8xNys0C4ICqAwwvwt1PQnvOGtL4tgf9u2sGDLsgMjTIROzsWy1AA3Dy2mZ24ql6zks6
Wte9606BosedQegYmdaBA9YtJsbRvjWUMuUw1VKTc8Jvd6Bec3CXd0wwrjTuEE2QLTOLKuSGrtw4
2zvEiRAV3Jlp3hK5VxHhkonVyQ1YvjsNlUCCVYInfYTtaH+X4M/48VP5QTqKsqs+2ByRMoUOTXyX
zMImbiBkl+TcAARiOHlB/NxtMHjs7alDSmHtjbrVwVfPD0oBB1y8UXPbH8fqDWvAxeyZjzUWuu52
Rzqk5lLLQCVrvxW+LnUDqVW7UkSPc+/ghY03cpi37mcVoxTD8suu7ZJcSG3IuwWoMs/g7XFZixcZ
k9DjKTkMgM6e7fU45+GwVqc22PqLex/c4HJ52M0bdoHpTUPvn90h/CR6pRG6j6bUWSLgYfg74MMV
y8iudRJKfAkOsY/0DWEwAAnMQT9jAq6gWdtiN18LI672N97BG1IlXs/97CKQqgBpR9kMTZiqDZd0
pfgAqolbu9IPM9IEDbQymxNb/Fu43gsWkjBbrs4ys9iUa5YssUeK5/MBzyo4JkD0EsuRB3oKamZg
QgjA0SoSaBYNxGBSnMeqb0VHqYMwBOOpcX8yFqdsEANL+1u92toOQxvhp7ygDV8G6DwjbGxC2n1m
L5M2oGcZ30tVGjKNLk6fMbdURjVpjBedCkNjVq3NyxbHkuYLbA704CyPNt8QfAlKRJrOKJ6PgSAF
N9sowzmAMuxIQ1y/IVKmz4f/8BNsSOT7x7HGmeM8+k8Z2Z+E6+mM36kMpXbbai7Q9HXbDKtPIIz0
rq12ZqJ7pecfg8ARWRS/yDkeF8fGnztJOkaLAEeOvshFQsK+rEezQLL42hMgnCLxULpvAdSmjYFJ
+YsT/6dulPZWs05dGx2DEuReIs3nfue9T30FrNKZHHhjkCtaB++j7hhp/Afy05/MH1iV1eCyNKZ1
+g5aMcHFqGWm7mLAjH/Gzp4bg6P/27kT2g9ntPlWZI1XgAUtlUrefmVjodP2vkyTWGigZ48V4cUs
6qBHDhV88TmcN3zc/0+sPVcZCLR4IVj3FJ3SlTlNxRu5qZpF+f9/xhWXZZeQJBXVEAiWeLJ5m9cc
34V680LlVS8KV0oo21IkBocjIccHLZp4hgb+CeCN5lNp0PrRRsm7QssSHJ/NGgg4TkkVMuhVSfgn
KuqsdgUcrWMw7eN6y880FFU6rXi71bfvtYfYakJnTgmrJhitZGLlccCRYdk4gSb9H4IbRCtAHzhl
Fe3HB7brsaqpBBR3w6HIgc3XOkAiX37w2mmZNbHXOMG1kIMIzfy1ZwXcnDoQK4qnMTfCoQFONqw7
dvuMB35wnzqR7ax9RhVgq7u02tsQc0VxszEEbze4dK/bZCgPyhKhPR7b7lxsoHkV2VMDKfj0gJKL
MvD6Yr5hSp0IgknKLpTICiKbO48Jw0e73JaJGBj1NSU92Yv0hnvBbR2EvI6VxY/tEaC7IojEaWsA
a61ik5C1r/1SZTtpsoHsCNIfxMc41jawR5X48RNBfYaiyoVvX/gndUcCTsB6Jz7bajkT6/mIZpbi
sAu+Gud4smEVX7fEyw7qhEzmamMzbJwxYkhbsUuJ/XKZf6rAei0+WssEN2mWPkyhHsbv3F6IsJAX
7GPwwXl56EvHV/zyBuH/kfczgnfmNKw/IHY/7t+Tf9jIFpV8zH5nMcTmvx0PPBx8/4S38H6dL7mQ
g97Zu28T9frABoEcpEyakxuojYSVDCXBRhGGEhSvbQax8ZSJSRwoPhVXBXJ6PlMga7RuEfO+mjLd
wZsi4Yli5+94NsqOIjh0e90r+6JiLYTDOAof8vvIFtYBt5ZhEcuJgeFQ9nqeIz+Ce1e8gfv902ai
A5kZNtIBYUctQfeZnPd/fnidDq1KRBkSMKnSs3xDN05xObpDU/rUeIUilphn1g6QYNPQxJwoN1yj
dTVu0Wr0P/OWn/9EnFbPrKFuGc00Y83cxFEuUltX76kzd3uaF9XepW+l6kjFUREGDwHN9cf3Ie9k
THRSybEsP7QNUES5TjzBTncbhku73ZiZYE8WZ68rItkWLWH/tJE/dC2To6+hSom+5L6NCQS/dX1W
1qNCcj3lnTmKzN1IiicVRqNQ6rYwEIu6gJpHdnb1Hy8EHqosJqEhwUgKznj1orZS2jMYBJxy3S5r
1bb5+6WAcz8IqFhPyTdQrSaytKF0bu/ezaQE62AAVP2z4uGntZyjO0P5DkvnMbNYJBVRZ6JIMgCk
RIx4MrHlKWGn/dGkNC5aqBPr/6T1ZVUlqcjzY8Nat87dGse/qHTPSpXgN+Qb92PxzQuo2/Jkhvib
bzjV0bb+w/GBHbysBa9ITLPAgV2q/LVfJ1uUyo+Q40yHnYvGoQt5TyFk5/AuDC5gag+z5bl4A5TW
AtG8zgbYlg32cvGH2PJvK55II63xp6CVAfKhXtqFRMOkLLgbrqlh4kaJPxMxNilibT1j3mL3QFtx
cBEVAiesojS2LJN/Cmpxado1HgP13lk0JDJhOowSkgfzPRyeMIVavC0OXNsHn5HxgwGFsehTIh4R
Y4S37X2EuRqfkDEtUILrlcZk2k8OjlbVhykyy3+Qp7nIYLFHZ7t9RwXQRJTWp5mYO/N6hdvDz/uD
MmHLsqB0Wip0Uob9b+dch9jqmpYeDoTQP219fT6eFKDCfIrDbX9saGiSH2KSCdL0N7AFHjb+4Vf6
bzuaPIu6KqI6wwuC07llO+ovgQ3La+CcH0Nc6BggwKAMxtIECEB0IWuT+ozlQ6CqAkBq8lTEpD7O
X3e0MSN7ML9KL1rs1+0womc+ts4wRtxjbeWE/NKGusMB+i0jNDepF0P84NfgmFoN8QaftXJz5mbN
Co7uhQvLoHBvOEpu29c6x9ra044KQ6ZNddDrsfMfEN4HsWTZAckFUmi3TRy+h1GKghCameIQ2prm
jMlq++brQonkOD9XFpC9axi5vIvR4QHKeFfMdpGPd9lW2kFK0u+Kimf1IdG7OvHSm8s9CCSMkUT7
ft1doOWnGdzBqmRN/zNGWWzMTAr8RoAt8D1bXjP20p2eJbhmjhyAWEMPK2OUpvSIVihQaZ5puCVh
HgcdMww09+utKuzV1LsUpdFj499KdxX7aHFbl5Nyr+SRdQjQ9XQn0K52zE5XB4GtTaxt86vEJZpI
hnQT4aXzg6IpFjUQL3XMfZwF5MzGfTwFriC2+fEe9h8H8y15evILKsBXI66u9Z7eN/0lriFftC7e
lbynxKQNX4Ab6TKY6mIpC+ETKKuR0iKX1yRpzhJlfazTseUx8vIL8lU/1+m/j11S3JNhW3LKrASx
ZF6vUQGxh6ivPsEA3XK170wdhwbYMxGGKYTq8VBw0VB94INL/oc6JAnUd9dADQDE+ZdBjdX6OIZn
HAom8w8PnyvqWtHRq7cZWBrfCq8DJfYtCnPfLCakHIKdmlujuMSzJdijKHCYi5MG9aA2T3/xgZsg
MCKZFz4SJ2SbBNpv2zljch85I0Y1xLXGD4Ysi3oYk2eg4Nw10jIhYmGYBWeyFtnq5zwcE4ooD+fT
9Y/hFKKeYX7pjpGzEudmvXStBTxuxhbfIQETqGzcnLaHJVrb8/3cOqzRv2ZcCpbxMPt1lwo8xQxB
XesfOG1w7qOBA41uAIF4+5k2y2BcxtCeCQ9IoUH091cS3ef6jG2yOmusMmbTjwPvDd7fDW17310b
1oNPgXYPYbuMNnhkJ1oIfSizwtxoYDzVoTDcwCsI0Q1vsLym32uCtVe1CCzVT28wDLhp7ZS71MYf
3mfTeu+Misbbs9nuupALAJ1nxdVDOplqguYrGLClOAl8touyA3xLxeA/n6L1bVicfHOJ1jFjY+9B
j2M/CkAs+ByH+toiMQ9iy8QGA2+K5Lnt8ZTablf3KrC9I6AqpaOdHvb/jAqGCz3YnIpgmqRcZBOt
EpDeYf2cmw/XVeEyk4AoxjNp7X5zGCwTykMQjTYJqusEkxbfOQEtuQNj0Wl7L/E0PVEeczalRakP
sVgCZCjGMDhyMOzyOi/zej26h+MXC6rDo4WAjy8NcMNSiEHC3sBZve5EFmTmmdBkgjWjm3myqfEL
uYY3rYIDlwDtw4dOcPLtuDM1PTcG7E7+0+sVaEWn7SVBbLtw+LhnjoJGzZQyHykD8pZT1vPY9mfQ
WdBJB9WOh+NKsfy7sJ7GYwUbMbCr6lQdMAsGlXibGkvn7lwYyQj1kTDtS2fAlcoHzVb0YyYqZqaM
qjPAJaEjoKTZvhwyOO28pSwRWSrNV0Lqz0YZQzGH6+y/pzG57ul0O+QAyAzdYugcE9uXH9f6Oikj
e0aN6dZS1Wx5OomU3UzCdSvf8/tBQViNEbcrOfdBDySWpgxoXtT7pondOFQmq2SSF9d5Ay96FEoW
9D/3Qv8MIWh6SUJNpXvAHwBkqdkdTMlhDdyaM+OaTJpuYRaGicXj60dCnGKDXaGSTPWGLXxaYS2x
2+q/eyxl0/sBiyj79ymptFML6RfurERhN4Lk0DNlhdOz3gJpJTrdSytDBu/o0w7f5+KJDgbJfTYr
+ffZsFX7QQ+ktSoNbB6yIMYFK9LMJscsx2ACQmI0zbqdbXskOc4hDD9ivUTzQBjXP9UvY3qHlFQm
sAeISKVU9p+EzuIBVnFaWkw1FwQPbJ4jpjFCnufV1Cb4PZBJAXfNn5DwhXU3H/hn3Ackx+DnEKSp
fszNeOEPBmqy8eLcYPfWVsruJW5tQSTjIYgjRHTX3u2uQnTpEYjLGuViVPe10YG5Pkg2Z002JyK3
NkTUQ11Pr+A2k8aeBr1CBwt0XZc65pDkSoTIrQmHN5Ym7SPGPe+cmwl7ov9yQccW9CS+fSwLFGWN
C5NQxldPJaLjTbvZljg1k8hlMbKQq1KPlgw8JTOi/+4uzdLWySqh3rnuuxNzwgVHA8FGNNOl3bzy
sHhDfFH53tLl4/g1riEqzga5eDANCwfII4gQuOro7Pyw9Aweo0KuN8+oEgBM8q4EiXLg7y2jRAvT
7jJ07jhzLCAzg3RiSCDir5tYbbkn1/+fBVSkhMI4cxgMaeHOvO6byMGXuwHu1yjLJ5fEmlNNPO+j
Zu8fxfpWVRNwHAOgaN4g0XM4QIyU5YNdGIn+S0eh5jsFwBsJubiF0xEgZvIftIubbK9JCYdqbxqS
WZbISk/1f5ajmv2RtbxBo/Thz5We82QzZtdhe2kqINAe14IVV6H4BqXTTehg3Fm3ncDQUSWAi4jo
e1ZPljQlDkk4YYfL2LVvhPr/LmnCddaQrSZ4vd2KLbHzoTl7zPiDUdPJtGh5Ch2dQh655ti8fFmC
gF0x5sMqlZ7cYLtVYBvhthksxo2hne+bVBr5+Hws/pwqbjkEL4zbaUHM9Q4h5AhGrzR4lymH3UIX
xQG3Eu+BDaTRsKTeYdehLxM3AkmaD5hfBB6q8M8b9hklqiFZymsbIujna+nOGK4aeDE+55hKufLA
svGExIkY3M+q2kFTa9hw+fv8tiBjG4Yz3qWAzLdstXztN44cQ8hWXJDru+iP5xpKCjNuNkZXo01B
FWH/OpWg8UmWZazdDm24fdDks3c42NhP+Po3yuTfKjaSfoNi8co6x0eEoBphE97SWip5zL5q7/zU
01mWuSfiwc6dRDQCVAHiwme9KRmjcZPj9zWRYdib6tveleDznjo2W+OA4CjtDsSNTtLPFDua1HMU
nyh6EWEUxWeguHH+O5l/xIpVoKVXQEPu6npEMkGJFshx2JM0GEBm9bwBSNVGdp3jH0GLAp76Gys9
wa3HKQaBNv8JTZFhBwxROakqIyDkJx1oayqjflR9Vg+ciTHDa7L8b4T+/lxnG3lEbHWdnSZmcR3o
VnOavjAz1d1xP8+5tazlGIMgkOKepdZk65RBlEgwvFseWnhMrC+llhGja4lTP7DNXn04Hbljqa/F
mx/4BfuDDh/ZWj0GUhXbL1prq8erJGIDiiR/1CD9Yg/yH1E1CPIq0PimQ3v96rO4+TIRuNo2GnE4
mIImISESZMLQkUBzokygENnN1MPe+qtf36xcngtLCFzSDw0Y/HdYR0rpIRPRDzp/ro2GBqtzKhHj
z35ukl4Ky7DahVeQtbCIL7XS2WaFeHq5VX+I7YoOLdT9LKT0L4P5KrPsm7dcLBB9I/3I7AiNUBs5
97v654FHf+q1WNySKYZ+dI6EAeHQnAEjxKhz6PD/fUfbM9EXV4TLmoVB2ahIRfQWTwQLwIMeCMnQ
mlcL+4/7kSJ6T6Jkom5+OeAXMmrZPJ/7T27WrEHZ5qD37YRZW8YX3ZJxsLcuWG15gdzsfbvAhGd2
TgB4FqFuP+Za6ZuNZnT85vvZrXQKcyv0i/XkJdfuCVX69773t/uvOWhpI6g3P2zdCIipUhb2OTKB
uwxsAs9VLk2GySLMYTM4RBLBoawV6djU3tMtZrsFAc0ihiq/9FjidlmjDk7br4SEDHR59+zxcWlT
uUjM+FL32Lg/ZAYAY5oKA0Adtrr2vaDlR25vEwD5Ky1suGEjGCnw0DpWPldhaJwy0cq2xAuUMYAk
aHDheBtWOdwXPzDdnYIDx5xgmKsJCzIBdj4o+rx6ilZSmknbrk4UQg4eYqH4wwXwfTKCy7Fjuan/
2OwHZWHqAf6aeVCmkts2Y6a56DrYxaepJXeO1VJiAYNT8SN9uk7KWMhRu5XANpJ46hNDTfID3ekU
4hspuJ7PkjjEzPcgEjTz5TbkN7iEs5B2r4RE0EKZkk2pBILMwLZoTyXOGIUymAKCDuIe52IAUYlI
hItyO2j3bSgoKwRRRR+5zlz682JjawrbpaIn1Zj8Vgvxfji0HmPsYYd7DAMKKCvuPSfs4p8pfRxv
5cXkqHgEeRk0i/R41A0SRPvS1DqOSddSQfbhChEMCEnOMcYPKvZcYWYLJ7Cv7zyMpTpZbI3diV0H
bPDaeVyEuSe0RL0xdlYJjvchZyBG9g+3COwFZ9BH+t2bRjGa1ceTXQplsoMugDJMRThFdgtQouyZ
DDW8OJG3g4Gwg8vzgs4TBBXIIzENxXDTMUJ24hqWcyDpM29bo1Hnjjqg1Xdm0Tij3uKKmu6KBp6s
yN7cZ+16AZu/X58kPzMA23u0S+XrRp0SNjxwykECRs+JwmZH3MaO1842Z/J0TQO6P00p1C+1QI8v
lIOiVNI+ii05e8jKB0e/BU/XPafZJ+JtgZz5Sj13OYYO16RcA3HTKTMgQaCs2b9bnHO71O537n9E
8xH4Fbxe80JYz4EJ+CcMv2GPh3nSp6o75Ph3OQ10o/Wuj8Ck3YPVIOxywhsj5p5plLjI4UYvgkGf
zpUCE7N6au1VoTAd080bnt5S2BKhwaPC67ld4FhehZTkFQKPDxNwgTVy3+jBAjK4UN4wHagJO1fc
eM2ggN/iCaGCWIf4QMIRfr4rGmrrw7/TOpkKw+mJ6gQODYadiwqnjcTCosmSfJq1cVNKvLYsUA2F
q6Ci6lqLbpkruXE3cBdJqmKjzCzw9yHFZxFXpTDMsJaMOXfjEYoWQSr8wTvNyPsHu0E3mi80jYL3
hCH4VPcJaOZ6QOWpGCrYNbpumo99aXYRbYUKz/lVE41+OOX63Ri1KO4CSnO6lVpZ+Bdgd+IzFhvl
vf8qa64gqr92x6E88G5nPtayK5KD9wWta0bQT1BJxKgQMWoM7h8MYPJEAgyyEcotdg3qSSj1vb8J
KUq5rMb1atMkPW9X/kGaUw3uDbNd0UvS/eNHIMsXnbQfdOWfFEA9f6KozLwA24T4A8iCibEDg2Xg
JJfKu7i3eR6YrXZFhvXxXGQPG5ImppFJyngBwcGRTlDQ5WEvZBPHJwhwazNftleBWEgJp/dMEXCA
vg8ByC+v+pJrW8Vmmh6FmI5BUBfN77ahtnRh0Jg0C9YEPTb5+nEDMW0vhaD3Q+NFpZfF4kzQVE+k
slDZI7vU7bOaBZFjt91yfncT7fn53TJMsU5jYBFmScW5BNh2M7TgwkcgT7X9Zfs0A3gEiPhD7HHq
GLuxplUX+NwRiiAeXZLPkvLGB9xRppdrQeEi5FcbPB4yvVDJKOFppG/7QJ9Vq8o/y1bfArRg+Qgv
HzKr7IHhz/oBEziOY/q/ISlgdGxcvqctUSYNwfxxwj6/JQRpfkbxmfZxOhyN9jyxqhAZzqwBbWht
OKHho7bhB1lvaFmJmYBi/2evM862QggooIrB08yzR+zbaB19qGAdCG1zCHr4Ks0mXxgBltJh46RG
478anYvlFQIwyiLqdrOHw5s4Jgi1P8vSlKXiKpmEqxz031bY+jvmD/FZSBhTVY89bi54UVv68Im+
MJWkyA2rakMWbwbBsJD8XfVsYnAMSNThmOJCAb0xOSS8uNyW1RS+ilI9pDE9AFI/JjtpmWem7XIu
ZghQB1gvStv3tAFo5nScV1Oe7I1EwH9qq1htp+JhiODt4ldBbVkP8RCJS6SonywkXKsDvfQ9n0gY
gf2SPO/r5lEM+od+Hq/oP3ZXC/M/HxJinJM7eE0JgAtqJ/yVJFCtuDtqaJYTLhcBNP2DSHyGDvzs
DHwsx+mn02Je/Tcwde1iq+Ep7oJib85IE0w8x8jOjH6nDjrmcLNZhMpuugaRvT90UnsI3EaDYF13
spwwHh750aGJKCCPwAfiKN7q/gsOuZBvOxBRmSu1uZtxsBWOq/rKOIoXiqC2YzKpPW0MiP8qB0zI
7Cc407fGq00BVFe1T9HlFWNGMbgtlvOQKDQaFjkNW2P2TzE8tdocjjwB8QE7IDFcqO8DUl3zco4G
L04JoclrjjdN1zL1DaMgl+ZGDBYzEzYfIk+d+Ue3PAEFl26UBVP+VyxYxylbXdaGr8dJq+gkWDUz
QTSeD1OmKsxMxVetJjNpO5W/vY2FspOrJWVMRCUEQErQzOdYTN+DiFye49MoFIj5ww671jGBFicO
WG1HrbdiS3KFvvRU2lyTQ/PFGLWH1W9+lLk6sWX7LGn1JsG+cgWlTGmXkrA0Muh+AdFfTUXMu1nI
Zy3iKumyqWzPeXiR8tGmLL5DlNpuosYdxsE2UJnWWhPS7O9pOd9ar45kfRZjOKRYUpLo5djAVDy1
jiVXPpG4KJWucqqRn4aFpTFqWefhIfj318vwctavDJ2u5DKfybDz4Qg+ztdQAtmt+BvPtvWS+o52
NBjfvLUcRSkNMUp3xs8RzQQ8+NLkKYc3QMF3JASac/brKEnK8trlhMlJYKSGljZrCOXzUH9Tgxby
+bi1eR5YWq6UAUd4DhYHj+Cb+CXMd+nG0B2yY15NwnZUZM5YuwBv8CUdcBnWlO3kwQP+LiFca36t
alr6sMq3o/YJ3qbM53LnO8/aue+PvqUQ+rxpmJx9lWnf5XfjutXzIlKghPCpN7Xqi+YauPVn0J43
CbzkoTt/T8nyeWqCW6KiT8GRCAHA3k3BiXHh7hp7ALAMG+2BF8gF0gxee4N6SfrosUyXvYyJbLyF
q3tD3ouRfQADCixGR3ZjCIt8P8oTkoVPVCu4bC860J39O8kRynInDTJb6N9uMtyjqYaqvY4nyzpX
oktldjViZuFSzRIEkH1/72pMqltelkMltD78DXIMcQG//8/XWcgSfPimJhRKuwO51IlXb0SiV965
SOSy4Mugkv6Y52ENwyotsAkjjCWf2jW+TuMUGMgcTyomEzop99htqxMn9cII5V3h77xLsTbcv0lF
6ZXHf26rR/C/rk7ftuLNSH3YTuGHUTa098dVOf2VJut1iuvszRldQqnuCerK6aKkrAx13belg4vy
0GTxCFNun31i0v0+x8bxdINvnUa0cw1caqXeyYcZfUaf2jNTc4DncyQFEqEb98YKkFYzJ2zDolV5
G+6cpuSToNgRRBs1Zzy8rDhMfb0g4559jCcm9VhLYJaMxhB1daempETagw3xvDhlmVaQPdacF1Va
VaRpLzmHGiOVyUivAoh3vefvbEd1xv02LQhOngM4HxH7LdTcJDi0z3VI+eKFmVDErD9LV7BtKISO
//uCxzEBydpUCeIAPt6ccrVv3UMab5s0LU27KMXwGMU14y7SvkiGcy0+QDSuX3Moavq2QfxY3eJC
E4A7liq+xTMpUPGbyNJ7CmqvJ6sg2zPxK7NaIkO9gUAkDJU2NjDN90WfMiAR45aeTScwkEfTI47D
Hl389RMqOKEL/venRiV/xHMOjR9Fakh+i2PAaGjIqjEdwb9yjM/YbFiovE57sxko0HOHibGPzZqc
05hOzY/yPhiJSaO19g+AnrNJw94cc4sk6QJ1t2dGGh0zsZrlx9uoyouNszLjDB2SxDz6tL/lyq+G
8weHgO9TXZx82pz673jzwJQlm6Lw6PRa4XEVHjQQl8Rj7VElXNFCV2ep8w7zrOeOBMEo1z/FkO5C
dN8PXjDVaW4VZibydEMzPJb+WK8Hvnfo7H3YQxLaNV2LtExAuj0AXbiiclrDs0OQgv89sKKVOpjq
zhF0LdFc0ocj0K1lpt3yxc12zWYK+SgVt5HaFwLauFZFCuA2xQtdmmpgcXILMg/RoIXMT/QZBf6X
egFTRukbt63ija2miXj6DndTrLcQFuc5l+6pGYfA1it7vTVbHYPNNqm4xUL5AV0olsIa+74n10Gv
kkc0Q16LzWgs2mOghS4piyrk9VeSShMOATLo7bZ8wN910sJAiOXaIQo5GL1I+O64O0LI75bs6IGw
j7Rge/5JaCWwrmiyUjmy0z5pEOXHe1h3pg+UhJ4t9a2iFX4fBk7BI93dnWTYPUttoT1wOxqqYE5W
PBSIeZWMxxIrRPAMGiUDfNaMDrV09cXL9igwfe1FooWJpARL4fR2QdwwGPoc62W9ivuRDfwmpeSA
bfpdjREOHfFr6XF2EMfVm5rngJu78ggvmGdbYXATAHqaffGbXsdEoUwMqCbDfh1nBbPgfJPDnCCb
xqQ8tM8IhTbmYHLYU1C6a2E1B1JJyajKw+UKEYQHgLMekNtW7g9XeI8O8GDBMzYOgtHKpW3Zy+7B
J9rn/cHbzqZAJc+90I3IYj1KkLoS2nLlISm66SFah7psSXt44w/mRlCpvGXD6r07DctzfTxyp22q
5f+WQAPe0nsv98x3VduY83scveHktZ5XEQ2+mS5c+Ik/KB+J3a8LlyGfj26tE2y9TwX4oJrBdtQU
q8RYzMS2irGVPnyLiebInYElpC751QBqZt1LzqN9qJRwlvBiiiaVUf4H2MJczqPERfZu7fHAQguc
Z9/AOj0dH1vAJN1WtomPgEDUH2opCd0aBYkSn06Y7NmLY5qqD6DJ6zilLe8TBBvWhwdxbqXjU7nY
Pl2kcRX+JbzGMaH6C5CYlNwGtPpdLRcZftvIcOdQiCGNoXfeBNxk7EXBG2xXP32YBj3wA0VPF7jx
ebLJTb5gZrGl75VsV7h36vLmczpJg49GOh1yN3dRChrZIZ6NxOXAheX+9x42Nky40ztJNV8M3ytS
B/rrS25kTXhFL6+7dGNk0eRwfwtvItMIuwAod3i7w/r5YwV7mnaAISNSamauWJmOSH6v8z0g2DXv
Mmyd+8ptaozp2j54/Uaqz9+2u1K9iRuM7rEWFEIZbqNRwoFmUPNSMkpe6jnZs4dldey0AZLh9nkb
tjdTFoiI03zSEdb/6wml2VeEMNr05zlqVEEWs+BCh0zsOS2NsxgzIMboPp5Qd3RJhcIheq/K3N7u
J/nGFVOQ+ReZ8kzzPdFYsp4BTYMIZ00AGVprdr1c8MO9zM0GUdGDGsRmEDkcHzM+qVwcbC2oF7Ge
dokD/aRTMJH190NJq2kwyHuVmjgis22k+VqGPIlyrL72kVDOPcZoMbFnliXLeQle0xUIKKDeDOqp
l5CXUdfv6EPrcuBdz3c2X2kxGFOAj+WBvI/apJWFuA1/wq2fXewFSly42XGqTD0NBprs+3C4n2O5
jXO9Id0oevwioH4UrznTyA+sd9oi5kfuNduPJ9m+mQah4s0w6CtMVz8hV4zC4BlaKru0Yrpk1LPd
0ZDXJOXFYd++Dyf3JsQtLGA8yf16qVFQDlYkgQ4CY8EzU2zoxtdLDP6W6bkB5mBLqmLQOMTudIZL
LijBISTam4o8D8DGFJPIGS9uIOkS3GxLylav+zjoTEIC/+lK1hNH37tSsVvp3J5t0ntgh5yw8bfg
mmyIiquGj24zcH3dZ018rAflgdQRipYHisRLEDXjdMn7iQAhBQIdsrR0DJn9YIBjzJnkL31NEWUG
EhY1hkcxU1nzMRKe7LAQ0JoOB30ka03v7F9UDHXUKbEdFplm+rPm8UUf60+Au6YrckMuspTytRTp
UfW7QI6fggD13Afo32Yy47/mGV0FXfNFJrX9u/9rICWB+oYqgopcKVw5sdOTxH9hjbr/xuKREM7L
0qEHh+FHPUDMehXtWurF03cy5EepBFg9WjlA3m2b2UC97wqNcjdqvXQf/ewUMiDmpmeimdUCliwn
bMjhXmfxDSlE88ulwsZ6/XoAThATNb9RXdJI2N/j3Garmdg4x0mRVAfvxgrBlgjuOF57CB2DCsZN
gAK7Wq+KLgZd6tc6QhCkkQ69GuNHeP1I/bDF/4iNICqbypj1LkjR6NY3HLfBmpWKJHAy0aXzFgp2
eqCuBr2sxX3agIHH0Ex2ym7oZNBmT7n50soQ6+yM0uY69W1dtA4kVpGkwK4VzR/vcu7qqo+csh04
fjniKD83U0b6m2rBPpZMG1Trcwiu3tJxqAsozknsytgimMfmUxRBaPI19rdXGesXPQB7dB5GTTeQ
cMHeQQ1r2behnLE4d6D5AxYyZg+rxLkpQcAqH2DHvJ9AFJ+lD7bFh0v+/aHAebAH/GjJyi9FU4GV
rpALGunQfGQiXGlt/I7n2ouAx21FO0Jq/muA5b7Sem5qPmQW6xpzdWKlbypq6rp2FOn6ZfdN+NmQ
544CpdmCEUWOFVGaS9iWBleur4pFQjTi3ezAg+4H20RygRDasZGn4GeB8tkbHC0TrHUqh3UysFBx
Zz0OzRVtj7uDQ+0bm9ThYo3R6/CjDNQr8r4uyprdY0+CG/MFkepkhmKqD8LaIwshzvzBjbGUuxML
7AxVLCXiLFXCOpwWtAVf6VBlFKgAlgeyDBlMhln0EO2XXb74eizW+GpaNQKepOgXACIqnl+fQgTe
Hx6UHcIYbr+IANTbUGH1UKubNN+ckdNsdWgD0kDGbCATqv5ZFbCJ532hRCBPXWShTQNpEdJRCkIx
TvPmwhPXVcCvHdYPyXYXifMZ8iG/PDV7TJJReVc0dhfFP1JoW08oNNmnFcRvLEAHcIp4jITvYIxg
tcXaT3TQVZ2mvLwDjSfdNPy5hP9XxuYJ+6aRZzGYjcaTEVj6jYiU+38yXR5cVru+f1icVB+m6BDZ
bbOyBN6FR00/I4iAss3jbAYhlGaM4D751cS9d8K040KmEjWswLDLBqq0eKd1Avk9ZS9ona4jcMwv
yishLHsMZUXrlLQ4dfWoffVWr5F8fuIALkMSMaPN8ULIO/sTyNxIJ2Y52fXYIm+bbuXGrAQ7BYic
msWBWzI0JvArHPkgITbl4zGqWL+RCPBz1fRAW++8VNO5IU+NSd3Lkuxj6bGyU2M6cKuQsg1q149g
DjUl9Zv7AGQ2tldGREYCAFzDgRoO+ayBl31x4WkEtLCuVKYy3gpN34gKYzJfboeeJacCNKm6BlRD
ZD70RswmtLdcmegceCiLtNkWo68TRQP7fWRyFTTuc/zr88GpjjoGJ7/dgN0kAKE0ZTz/nv8qJ0er
32y6we7z281Shb808dKDW0eeeOyaNLkKD+ZHf8xTy67k5J9oJiXgjqQbf6hGk0QYHzITD8l+ydql
XYjGbBUvYA2aGpMEERUl8ywaUSqp51YUAyfPWihvvZRjKf9EsDhaqg+OqR7n0nw6NTsZoSk2sU+L
zSCjgSklgnUKvWpGZX3tzilZRO8HNQkmKxhw1ZNeQWNv8FaBdhohOgitIsT4MLxBAL4AFwXmUMC4
wGwtkpys+0CvV8cqvNz2DR8mlKPLnmRMkQX4fcibRZpCNSBYJwvdgI+ApDpCAKo34Nxkvq6jbVuC
m8CWX1TKQ2lZ2ZR/0NK2zHPJ5KWrePcp7flt/+7fETRXk2XUxudT5g7a+Yxs3AZNrvT+F47/h65h
oeylz3+PvdaGctRYSNjws3EmS1rfRYqNlqGjIhz0wsccA9PXp1OpvnIYUlvfY0Bg45Hr2Tdlnuwj
+cL3CQJfHFz/YCnpHyggxYE5MHmNZjqobtwkqjikYXhuAymBos1tuTH68uBMR46T1YU44nsQSDO9
UKT3e0Wic+nA3vUaaK+CEYF5dfbE1KH5/5U8d1oqhqt8LGdRJopzvdpiOBvNhZOfXpEQNxTB6ono
rLOfmJpZum4cbsXYMUwKrxJe9NdVLokbjv5iZci+tG4RLR8rtlBoGany5k4DTE+zHUpF2PbtTtlm
2Pm9vM8LCb1pkZIvpCFcMB9OnJwfCoyTCP36MXKvNlaL+EBUJozcMwFym/F0qsIEwzXOpdNXIzo8
UhTslrZ7fcKlkPSn6Ntm/iBxqH7eJKi90F+1J2613CtP+4qbwkYAW5KzJ164kSegyYGXNhdwmp5S
2E+fZcUIWQ1sDs218YEQrMcC3kaHwkq2+hGT1fEgYN77s1yCRyeCoy80a2TR5Xn8D5+gD+2LjZCM
Xs8UFwYIo0QrLbqEKCWnrLoSELo2gee1Wpfz9ENCBkOjemYDg+C3rBt/UaIeN5gV9+XAPqIk5i25
XAzYu91nC/ehpKY5oIFisSdUEkHx4IjhAXhheBB/Sy0ceNApet7UJpXL4F82xLqrm0Xup0qUpDsI
kjSMEyjP8HexxQKHlUhrMjX1E7uMJW9Qdm6ZfXep48YIUTtEHVTGjA/SCOuGBQi9tNpWSyeqCjBW
DmOqT5znee8LB8NWsA2AIx8ytyudws25IvPCFdaxXR2d4ZlQ4mryJ87VCbPPbXAaMi8B+MMwzoQq
5SskPgm6kdu0NaYgdupgmohX9ROGUs7p+0WJ3kHqxV42qlfLBEj1hM0CsW6jauv4HJT2HPRMio9w
FIULNwPFS7SwSeD9aXTg9CEOxA+JkplnhAbvgTdtF/IvoKWuy1CyrG+Ok0r5yufOOdYw6Rl6CjGw
j+Tdm146k+ZRQ8jf4VORcjrm4jHdFEfSTr2g1J/RP2A6oM73sBU2Kxm23fXWRb4GeUhkjGqW/mFP
JJEofJPU5xmOBqOkzRMl0QAQCqFnpUD9F0/sE85KGcBxjb5mLisLErKeqXJfZGF+Q0celUtij28w
hI9GBltwPVLfO/J0UWAGkXB/i0Gox/RTnE3u0ihGHS9RIEnBU8eErWdrdAqIg3uuvqSdkg7FDkfk
tn/Agh0Jetx2bQuXGHvaMRzgmpnRMplzsN5toHMmJSgfowmlLKPgITCDpkCl1c/I4GPBBj7Tgc/B
jg2h/+7bnvV6UgU/Z/x2AXm/y7hsx9I2b/hj+pG1mfs5cRe0r9AWiVu8u9brw8wV4c0/EAPXuk5T
Idjdd7WUIluy9Q6QVWLotSQVa5aflUtrfPfqyVIFCRwK0rAZCA9BuoLNW0XFfsU3kor88xsgVbE1
aT2nDb1vDr74YctcIC6yhHsdT9kITlFxTNmZnH1h2XmBlz5rMz3o/2oWW7FDzwbUqAhq9K6Mt41Q
uKrx62FhChqVTWz2KsQoKLw9cbseKKyzyj5/sKPn8qXBRD5Oqu/Nh5uf+T7WhS41jhjQAsAQVVIS
wv0YUgZGQQyueHjVN4JTWua36YljUTVXI1t6Pf2N+hfpGcFvY39mPElQ5b3QoOlcHXyPVs2oJb/R
7M6AUziVrc1hOlpgKmXyxotaEvayPkCx+fJncjE20vl6vhYv1bQG4Tkj3ZqC6RacSlbdxdHT0mri
PDZwdY309pw4P3mAQmVp585G6ZlQMJE35OwMDPCaK3TLW782hkvFwOLpOIwAR2dyMscdx1PUAmGC
71ArCkGFNPwKVDeO+UTJSdEHKaW/2jVI04WB4Gb/aPYkSVJyRH72EGCQIdyEY9LWZN4zCLoTU4a7
AnzXp0y4R+nV/uVyFbvnCySinM9D5j/xkmjHHsBbsNQHHKfs3f64p0fWUFRusDq17WxKTODtAVfK
afezv/YtZisy4i7EuLNtq45W/PxEvpqO2tdpNqboEhE+PlqU7BVLP5hWlaruQ63Yq+uvCDQsPoTa
7WjQIEBBXs40c1EKswiGWim70wZCp+iUDVKJxu/blm6xiOpIn5QjnVsXHawnWTJE7Ez5Ycim2t2J
52mCfwdNOTrv3xse1+7tAhZM95BLLaTVwp3ptcSB6DThdM/S7N9oBbj3PabKBbjLT+qV0p3yhmAd
AJpyQj+qrMVCaTj1oQ186EJ/oS7YhC3mLUf65X5d7lZwNJa2voKI2ETG/+mM12A80zxWk8Rpg/le
+SpFZUVsLXF2lcGF1Ty7E8fcxyv4o0bM8iGegXrNraqPzLuLkrELC0X4iP4BL3Ge2pN76m0pTbe5
S4Lig91WqLSQzUZzNEoYdiXtd5MUiSFe+Dj2QX4zFbvoI/oREItDXAeS0TgkxlW0nKoP4SLGjtc9
vd8VIYFRMCJC8e40OfwfjxYlVYnjqqWWKZvYGc2/zfEWBbaENbvf1cgvb8sphD+T/nOB3liQp48R
ilA9y12tkkN1feADWHoGhok/QT+EW6e1Z3MiHIsgaZfWFMa4G8uipr2FNikykbDSlMW9hs4KD2Lv
BuGVza/ldzs19huf7fuNtkahKksCvPTCgrM7UIhWQqo95P0rFhdd6aK3nNLxqR3sWPGxdk8hDe7k
V5hXd5zbiPNce0eGK9a3cZuVOslCRTAdSfipO3u4LC692nlz73raqTEJP9RN/QbVX5ONN29beB3x
Ai7w74AdNIUVHj60is7dUP0seospEqElUeK+S2MKUZCoDm7LPZkqMGA6u97avIdRmPOX16SGG6FH
wUd1xZHc/oqqbMoONQA6lKt3q26TBhWwlETLYNSGnbi8568swvfCyAoiDKUXFurJijuaj+lHebca
MJKzTn4Ict9AL1gs0mYd5BSAAPEz+oSy8mWz+L/CBUmYOpkNBD18eAeeAl5mZiwnp2VfSTyN6RuB
p+PXetxDFqXIQJaO2Ys8KoyBeCOrNqQqA3pJrL3MVQTpbNrFQsxaSl7GKpD32Y0hO5S0niIIfxRP
fDPH9DqPq+tzVzrOA1sj/cvw8h+eeHE9vhkE/p3lf9UpMD3fizRrATdNycHD35G3SRIDRUKdY8Ov
mWzyVwarrRLWYx8XiO6C5aXGXeP8ZIKqk2GsSB1RtvVmRk2H4zP1XiUG0oRh4oDz5GtDrcSGDSCp
wtfz3TKZrT3De4dwqaOKkQ5NJLA/bCdnFXom/3M38Azb7DHAQHophs5PFA7/ew7D/s1E80I43HMK
8ppsHwrUhv4rn45uOD/IGdRAhaRmg0aLqH0K//TupqcibKuRFwKb0FIzUAhz97aVh3HgS/Lk0SH2
nB6LNHdtnF27sdUB7XfJ6urJ0Z31b0DYF6q5GOzV2+Njc/CVnU+gYZoRZSEw3U8ideEbxhDpuCEJ
MRdSwON0dd9mTEV2u38YpQndcXwJm1ALNMPemIBbHsjORncd4OpKZnUVk4lWnAOAu5Kz/CylDc6Y
u/ygTENrRILI1LI67KLDX6ahwu9IsS9fRKEERl8A2Ji9+Lxj78uiGfTYOmobPXyFafgj4gs6cjpm
el0KBZcYpG3QwWYdOzxy2TXDW++/Pj2bEJnZZbfWfj1yQ92gPEUPzWb/DCiZMFq0+qB+8B45xofP
pIQv3RFu4vXMEm8VJglstNgiJb5GfpGilfM9IRdNYUjLpvcDPZ7xS8o1bwNnk2QItJoCUr0uQctR
Q5NrH4m/wancJQU8/gXEaruaqsPIiKfQY1q2BXz57CfKSzbG+nC5Rlep45xaFlgl8h4w/hROHHXX
49LsVDRDDHaj2UiJwb2KVd8flgJKbtl8wjdVd0Bt2VshK3kQ8m1d+lxDSwoFrmyR5sBbl7ujqwaO
ZlwXEe7Mk5ZIf5igf2aRomzH5lvgVUXReLiUdouaKRXe8iQkbSVma9KTVHWkuwfTYuaYr3bHl3YI
oWilt+ag1XyEixXbPjZwcVm3NWsXwJIZBF1uyFXsX5ZpwfRH7AolKzQDSFGmYg7HPC74fYJau9m7
5Bum/XFhRexvL0DBsJimsOMTT2LH2erHOpc29ZcmAjSO4AgRAf35YQHWoZHqZJTp/WPUU6a6bxCU
Bex6JTnZmpO9DMP+FUW9D8aAwXwlNiqwdMx4WAvzcUxsFrLohDtj+L/2lxAZux2gI9aodsATgggA
aFeHlWjeZRJtdON8CYXjBeDT+oswnQt4SHMJ3W40r/d+9H7d1yFKy1snD+E2H5onFqOkivmDuWeP
bBsy1c9qZnuVTU+OkME9cFW5Nk+/wCmckzBctlkWYh/8X2qzqpqA9uX2g6L47AVvJ8b29vwO0F1+
sbot0DuzlU1RCHvm1LN/2TbqBejOaIN+pftePuv8rKh9M6NHkk3kcBzmf0tBeWPfNWrLxjCjh6HM
4a6s9k15BlaBBZvMuRetJGlaJjjKpBDIExakppjhOYm/PLPajoJmIZhtWM+Vfl0CNfs1voVoWU8g
nD0FYiiYBpeSJOnnvBKUDrgNOnrWgpBUrKjdl8h292mRZIz6/vX1Jr7FU5hUjf/zjL3tsgfJNdNU
kdVzsxrMQHgp0zjhIaHfYU9v22xlbvlL28cM8IZcJd5Pd6PEzxf0AFpgvZr/rrnBsLbiazOBCy3F
asDFdBeJZQbeaV1sZVEJMpDyg+Y3d6H2E03gxs+BJ7bpoDZxvw/SNln+RrZQTbXiFKTpocOw3flX
Ab7ryAfcC4ncrntIqXreAY0jQvTH/M6M3ThY+EC2iQ/XzGTD08Ei0nVs+Cy5Ddvgd7toRZzWhFvl
vbhKX7rGrgdMHWevZmxqX/q2cFMniKrPwSgygrt4ICDfYv8NP9ZRMa7lxBFQ5zO7VHN1J0oIH9gq
PjEKXDXr9a980gGxsHIeRnDB3e1tYKnwi8HJE2QKS/2y4+aa6A8WN4+LJQ8vggE6s+3MiswhC9oG
nLXW0aU1rkFB1DKZHRNsU9JIdKQRp5wK8oFEfIauZ8WzGg3kWyDY3/zbvL5lmS7xVbJ2lB4pocii
o3XgpQxafkbc/5htDO5fGrw/Ngf/G3bVPtsN59WSGVnQlHy277fBPG7JkkLvHfOjsAoJaHAB+Rbn
3WUsyp5suq2cJiT+wQaZv83gLaiUfqrQ2/ee9/26WMpHvMef9ytxAEsaprhF8huJJLvgkIrCrkIA
BmnKMbhp5v9r8GDOwkzcm0dbjTTXyDp0yOjfTZTtS5wHmQ15fzPA9FIPVJGNz25e/5v3xNDDe/Fp
h6zftkX3DVvIbwUxXlEzlrFxOeu+4pg7Al4sugU4enGscEHB/RP7ErHwaE1jyWWPUz1YVCU0l7nL
3TgY7z6eid/mPsxSaLUZdv/9/pQOxs235T9Wq+j0pmC1JuAYTgmEiiomGOv+ueIL4r/gDvmxdIZo
PzxR+17Ceu1pCA7GMoxBx1uXR/wPRYVjDZhU3PC9/lsinaaklc+R5zvZ6H6ls68JGRVTFOTIOAlW
+J4Aa1wqXIe3i1T+kwUal1v76epzq2pZzMW5OgO5themgz4OaU4/+fObyzwlSxvV7erq/POoL9k8
XOZgODbCRLfkBwU+P1y4RnfZm5lcFNCSNnJbld3jQRlw7YTxVq6BaT+tZ9eHAuIpsmdVuvspjgDZ
bqJr5K10CSOUnNr5Do6nCw3DNjR47LurnAeU3wXvb/JtZR21QYM8zw+x+k6MCWC+RJmH7QrPN+cR
AHoCXS8fD+g7tMpHY1M6fdVnZlH2Moem3Jrjv6xbwyIfpVBYEM6o3omO7trKZxvx5UpOFUEsytJG
89FcINpyAC8zCoX91l9HgTh6X7wtyvd68fSAWExFU6UPp99IAMg8zpVk2wl2F5sEaXlQOVRyuDFU
YeucrjMNEF8pHUeFmvF42qjK/7OEtLbYltRdpYLYOtGk0bX6S6zcLCMeJnkcCb9hOqX8f36v6U1q
qUwF2NsNHoChYW6287pCQc9SFYa32PEf6e/8i/FRJcPAmXLGrDI8y1H8qJTvr7F4BRIwwdBCWSI3
7+DaO+Y067Rhri/iquteUMzQTWj22wUgUiD3FZ1oqDqnZ9zIn95kPbEC90/HlGNb+cxikKEGqnuM
m6x5VEG1NKJh0oEf9JAPLAbFaSwG5XchrdOpqch7fBoAiam/t5vSXND9tZqJA9/U7i35wRU/bEiF
Z5v3YNkEYoF1tu0u22Tk6qVNNQnq2mFLKW3rEvAtKlYpw/kkeuv/Ygzb7/Nzj4h4Pg7/uEcY9/T5
ukK9HEW9Wsyxti6dX28RR93lqO88DXrOjswbd6tT9tFQQOV3HtCBqFPISMEYjXgMWawvatfmm0Qq
t/9cUFpMHHqcwganj4TzAb50avTZ0PXYPfb6N+FY/iT1mfLqY9+hRKzC3zhjs/NZ8hWLfnHwT3Aa
Swy7+cFtV+kaWMnv+mfOsz7/jPm+lbDPNw3Ib5MrPPRXKZiktZX8NwedCnDFDiFJBbAGus/+HpaW
+eG2j9UHCKXbB6Qya0TEWI4TV7RC8D+E5QoKxSg3jvnBgtrwd+RzMa3lw272Wn2969wFzh78wMPD
b9G3sNjEwn0GygLt95HZqFC+CQ9QnDuixziNp6SHGXb25pSZ53C2/lGlvkiUmJMNKxI8+7p+UuNA
MBbzwExWrq66N0te5B4XflkkZ+BMghHLA2wOcofCd4pJi2JrCw5pwHuUM30L3v5nQAD4BJ1AE1rf
SDW72YdQTMILxj3wYiZt+6X+VRBlKIK4HxBLvy6x+9FCNlG5CUU9VC/zqAlGYsrfU8SptzIRvH4E
6rkRrUG4EYiw+0IIQ+VRIUmxyS0IzgXjw1xT1Pu3ImWtYrHvf/Qn/R2am/B2UAo1ROdCaCRaVwJC
Pui+1E7liSIGlRjxRJ4hgIGu2K2tjDJAbIF4u/zIbFjQ8nZ+ddeHkvIdzzTZQQCxcwEqaiLhDuqh
gKSv1vGY/u/E4UuXbSyjm3WKu762vAhICN5hFKK/i6u0iL9ECd+O00RJZsoep8xVvIg665vR/u4O
xzzpiQfWPkZT2VJN3HZtO6BzLfMlvthvoesNFpCsYUT9HPEZzIeayq0Ze4yIMOMdLEJl+Xu3Kpso
2SMjBF3l0cq0N3bA94aAb5tQqniWI9Fz20ppWUiMWaTnY62SoUeRvJS6anped0tFs3me5mOuO/za
pmGYQbWY5OjaTQXndBBAvf4ggm11rkt/ZCULhPqZwAEcCgYQOYmepE+sAatcK8MaYZ5VxF3Tz8nG
YuQSgCIF1f1bYIKb845T9pVB9hx85tQspKO2KZ4db2Js+qv5jp9yo1EovxkWwhPC1lyDyBZ4fSAm
Kl3vQlCM93ESmLGWwnShA2/uqdBFWuagEJ8K9jWTLHj3Z0Nb7RKOwoQbJ0pdsl/0n8IvLSNL5MUu
zAyE/fGEnnu0lBInPVO4cow58vsL3Nk81FgmL6/ORQnRnXZgqzOC7LxvXTItEyYJRx6WyR8zyA8E
crIcstuGNiJA9lvHR5+M7XdEU4+BVijWxTNCvxg8sckU9QYUbGMkwLd4zf7N+Gi1XixnBjKCjMZW
iImwdx8YuHFkUFrqVvXswz5U66n9VcmoYGgl/epP3O2GTJ2iLF9Zne+VLIzmyeej1rxgUkGkiupU
8U/oWg8n/R+Q3gskWxrqENDu+nBe0OIPj6dnGG+F+zNsXoPdnDcK8XDJxLuurptvCa4BO6sEi1l4
IoM0SBuAbMMt2bQQz4WLnSyna1V817EpC0uSuCaJg+j6VsKCB+v0LJSh36bh3NtR8lyUf+CAkNdf
xd2HrAx1/TtsyG6gvc7H8NdJcGohntsE+Yp+WKoM4+ujRH2Qc7NIEgHWmiXbZopD0YCVBG3sOtsn
U1d8eqEnlw3KusynlwgJg0Uvuac/J/EYB5p+4+jlcLk7S8q9Xxat7N0zEuM4Asc1/Zp4Q7V9Mtbq
uavU21DUtYoUxzYRWKApMIjQGygqnk12L1v7+7yQTUby+DCoIPQvwHhSZ+m7SA4plZWgQ0782Fy5
tJV5Sm24R1DrVU0mUjCYTsa/LA1w2LmDd7NxsTdqaMi1LzK5T74f0EwHdXIS7rTghdzJhvuINoEw
u/9UhNO8HP3N2oNXUDDWrpWuEiMSFVHMMIfQh1pJLKNZbBF41TWclfS6Ov/WTouszZumAe31nWBq
Tc0ftwpMgeyuNtO/AU6c2QVFvl1L1DEqT3vkTr+wOh6g3ZySdHwO0QRoSDYv2K7pyh+tP0TivwkA
jloSdckwi4C4+ss+Q6Y/AR7Ov+hQ3wq93fZedvigYUK4/5RVLz/UBlA+jYzgC42puU7057iYaC3K
sivzfhnloFbBmZ5OmRDUYS2zkN3PP+UTJsqGfWIBgYjkgD76V91jXDh+Q9so67mUczFh2vyIwoWS
Z6N9il5wbzFFiHehGLgl4oXdjQWzlSlYd+uMkgma5MEP10u5O/T/9kF19cYrmFUG6e1iD55Fj7hC
ojYc38+TT1mxLv24JNuesbn1e30FK9JxzxUVV/WBDai2A54x4MsuejndAPncRH9C3qqfGu9IFHRY
VovAEU+gKelKNaIIPxypSvs8C2lAPQe3N3VeBbVHKLorCYvvkeqO72DBPIGKfivrUSZps25Pn23y
PYLcLe/euH6vf/KfE35IBLAZBVtB/z1FvcdMvJ7um1djhOBRtmOu8iQ1CaGOen0mzTxTk9sd5nEb
v6F90dqUOdWiiQsFVmlYrPlXgzRSjDRGpCZ+RFWEX6j+ZSqG7/NuPAjRJABpaaA+mcY5JslQNfFc
oSu5Uu4IwF2net3UiJyu2tiK1mDiMUUD26bmsIIhWoncJDOt0fMQAKfagw1qySv+xG42ToQjGsT1
HCoXDCbZnSvlg8A0W8xmMHihO3LNo17gUVrFV2xFeIvjGBvQFIQCMhqBNZ7pnxc6sG0QZIkLun4/
7lrDEWQi8mb6p6USnyd5VTsrT/P0NkfEKuNwkZnw5f5zP9jILOt7+Ki9Vj4+cnLsbD6vNZqO4nGC
60j8GEXGtr/JcxhUOnEvs6qQAe3d0tqdy5j/yR135S4BLiI15u/CeoQ9skkXvWsAdVVwDcxE9cT0
akertspHRAx8Ckv8ZbI0+ABqe82OHfbdPJnw7W7buR4zQ/iwfmIroaHQ7CuTSQ0COdtqyeYKi1Gh
kxNjQcrl8GWWEdV67/wIVCInd3UScIagGfueRZZ0+XnrbWWmBRio7Pc39+ezFkla3NDmB7PPrx99
1mAjOYwzFQrmRx4A7RyeALWRMiSs+ZSRDKMl59USqoub1cnXA6GfWhtQ1x+zCCLi47OeQ0wl5+eR
WnA7pg+eqHj033XWSNhOCUo9s4iATlpUHvxA9MXhx/BPAJvvCDHR3vocS8dIw61yWf8gzV8/BpYK
Qf7owfL8Mw9lL+uDocIYOTAoNQV2ir/QsMGlQNwGINK5Y0BP0EnA+t0spi2XipiNw6T2Une0yyTc
/SOmuvAQ8X9+B8DlA7Z5MMLEXaZiLx6yMgm2yV6yBgshFNnvY/XC2VLtE4d/a6aLVrTCqL0B4hRQ
Y4w8Qi/v+pOKDLNa1CPYYVtEHB5mCyXn73AkB0wSOmP52P9zGjbU3vfCdvBxIZCTEZYyubf2ua0e
ZyRC+a+MUFVlXbHDrGN1LzMpL2uu/g5qL3ZjnA86Z8tcdX1ERZWhSlwNxLQpfIIJCbZhBC58M/gH
eNN/etZTf1XMhrIjhApt4CtNEA3qJ3mPUK2r99EZM9uwOJn9E+EbxHS52/VtzCNIXHUCmZxXNuRm
4QDI+ELVMdO0ssCgEoB7pa3wX19BTm9fpcjiyot4Tlt+2/ymScGhfng2e7/AwcQbE5zSHC0rolPO
NsD1DM/BPaU3o/rJDnYahqV4ojdNufoWSodIPBBli+TX53uSYeFbOldq7EQHFM5A93fmIdThCD5m
J12cmfFS4bbDaM9SWg+gI3SREwV2O43I7GnxqCKgQs9RY0Z2uWuN1gZewhbhIzJeAXdBH1+ZKCY4
c9EDSxhWl5WeygpZfo06KxXQFARalkAL7EKES3PxFQevmc36IH+v3JgmpM4tWs3f9IHBq/TaGH5S
BwsdY2TV+cCwFPLzGNAOYp6hfoXdGQILHLn18Ox43ZSeEMiJzPTCwqAr0wiMx9ILyCT9xkE8CUu5
aieNfB2fTaTx6EP8vF/VfU+BXJV5selFt+/R9kn0Yex7FgCCE7iBDyw6jRXTlc7MfUTzKixAI0Gj
OACaXU2EsrLVxGGMxGhx89tQWwsz1+cR0ItZId+6QrWj47e9N4uBWL/QXBxN6Ddcsp6werAu0/GM
sc75SQEI7D6w+EEodrdHH4ae6JPgksiYwSLaAuNDvY2FIwV8n8RkKS3+aMIkJwX1ytKHDUuSeXAH
TOV34tEFhk9RJPBGuBe+t8Ps4FfymthFmgsagWdAUYVr18UUiGLlWHWBZeM1oJvjDavv8bUpwm7x
lHa2Xc4/Tsj3vW965RoGJZW8fk3sVj6IZbGnIlPVP8Q9FaWmtAPj8dyg6D9uj3lA8tI5JGiaQ60m
hJ3uXZ/3rGxLtueC5breCK1nRe+M0xXwLmopke8SO+WznP84ZCuqhSTBtby/pbOCwJIy1+3mp3mG
/l7mQavdYzMZmjSEhBTsx9XiRMXAgCBbSKQCPX8XcvnLRf7DtpBSn6gz6k/qNcfqAWec2B8rmCAj
9ZPwVyR3bOcGuwmH90P3Dnz9WYJ/fBj78rILfL1/FsZsfVjKqOerBBSNSwCrxxgNyC+FeGbm/DDC
q1j0a93vFEjqxlaFhYjmaMHFANShJJ4AIUqroYtImgaRzickUnfWabZ4UFco/67RUFrNtTpkJp8n
tnuL7R3WBMYdn8x4TQG2z9dZDJNCOCyF6irW0vuJmNtnbcy1qSVWYdJQ3wjEffxUVgaRa04uNCvY
D/JP34y9MCHO9s+ngNCLU1c8vQYFQOB9+WdfUTWdUOy1Rz2d47GKfG4xSsmn5sfxhXRVrpEIsaJD
qnpTwQAn3HPJdkT0WsvD7quqTmgF2FGGy6cvRY2nBtNGChCSNpQRNmclD0+mJs6f6N0oG86sA2wT
3S6hGPIlHNHWYT2VTNAYTjjY5PhVBum3b3nYrDzf1o6X0FxCclZ+c0/HM1K2NOlKnQ7QaEhXmYi2
bHsGWRePJ6GioZ5ADgeBUH3eivmsKitmskOyxLZdhgJ3uMkAG9T7YOeAiZQ4iwDd7YN3RT2GjRvH
vaJHMlLue446nI1St2gpYcFEiQQRtPTv3jfv+c82Pxlcv6QMWqnn3iEP31TZVy/ETHFIKLDvFMNc
K3O7lIA0Ofw7fnnLcppTRGvLXtShApRwZBWZyfw1j3rb8w/WjUn9ZC9jHtUz/DAFSMCC5CU/Ixe+
y42JYhQPAnAp46y6y0L8QA5tAQ/3+IxFFXMvTdQRjcp4olKfva04l6T851vPVdP6AQR72lO1Sd/c
qsyj9mGZCMpjhxiPoAf3LmOLLMM8S+KsNGKLLk+VQOyACWVxrVQVKrPGdD7CPpx9wlvNo24UXXga
/uB7KsD/AEg8dTPe1Jrp8HTVpcXUY0pOzHh0SEKHtl01SDNWF5qiQOjZyLurexz+6Ty3KbRRodxw
gUs7BnEOu+t84bsj0vlWBp1QTbEYhTtxOUf0J43OPh9mEB83ErMA5n8ewODM5sAVpzpKhmcT/Ti1
Vu5yhlGsXGAfXq3G7TlocGCyw8iJ974/VSQ23xyWpmZJFpCHHZf9UwQkMfUeCTEKLzAViGno7EEX
Ymkm+4HlEer5o8mkfrc7j/A0Fk1EwmgQBTBenvg+1RHnhNVGJd6nvm8Nq0ECyywEwgBCMhzmKeY0
PU4NAw3dvulnGB9bz/xwuHxPHrEjkGlqrd9P+HlBH793Aiv1vqWqXtYaB5bhfK1rNnK8L3K6iWVO
coz+GSnzEvOk3raeg4GKUVJot8qJhfPjS5bDKTqznjHs31KSeoodxAH1KflGeT7zkegc+U38yz6K
UEjyJJm5fhtBx/bdn79YDl+8jToBPcU6rdQf7DG/vAZ+SxmCqbMtk2js2bPVVtuhkK1bb+1Rcipq
QOShpNI9SUn15xcE7jIv6UhHGAJitL+h6wqcgvrZ+goLnWT5zZaQy/+ZNCfMUPavdkGds4nMd0tK
iFNWFLyprR5PwVJ8VDZSaHGuTNx788CLbWjwqBk9CD59KC/lQ43r7YaVD/D8TI4wHevnf/80EMOo
ZZEBahGuNa2v3JF8+O0dKFxP5Q0Die1/lVettvVaKbbf/h56OaZkxCUkXpafVeyU9VBS91Dx1tcX
MCFtYhNU/Ha0bGDiA2Wsg1SWOgXtYBnzSM+ZJtkC9rRsEhNzZ+0Nb3555vFsPYHfRgg17AxjCgiI
ytlTIb4ILzD7BFDwAGn1tfFJFo9dqTyd1OtCP4N1ePYnVavtrN9frXZXjiY4o0zs0aC5hjHbMURR
ttdhpQu/ReTwbW5OAtZPL6Lzd8/3zQHhdL9ZAM4RinUFGxLteplLWP2H1DPZtJBxc+AKxgYPTRWu
xQZR4jw7eqS6b63wDvwWsq0fV7akxhcdt8Xlz6iIVMIASO/ARyDZiMIJkX4fBPiKEMK0KybmrQAO
0WHUrAG/GZvXPGFPogvPZWyd9pwJ0+3hMeUXZUMw0tLo7r2Ov4s8uVgzWfUZVgnyWYJcgARWeZWL
wIdQK9+fetrRkLLGkgABRYiNNf+azEsBaX2MXvF8bFjM9woKp3YUUesVLRnGtDHHT7bcCKB5XZCa
JIJhtv6Lx0o/f+Y67wdW6SLtd9SnuCjB3IqVQri0RNnaJqpM/rv7s4x8bJXVP/LZdtBWl0dx22ZU
j7X/XmfJt+k0AZfVR5xiKyyX2L6hmrPIXIyoGtY5/rYB5fWRJseu1ND8PONUoY67NFbrwQPHWlmW
DQuBuVWQ4Iv1Tsu4xMhptAGtTsOVntLyyUWC7TBySFT5PTlvFf5f4Sowzct8+QjjzDwpKbDqWfbC
GhRWH/qLIdZVUY0PHJeWGas4zSiB/J2u5fNjJ1414YpUb7ZWc7vjEg/41ccPQ4OVWSVgMEeCJ+eR
S3piBwdcVLCjvIw0T/yX0deGnL82g3xIp4QttShB2ZFX5nf9lK8dMK35muwgWiipaK7eO1q5ZpfZ
lfiX2z4mYMv67APlOM0smVJv4d6/kQh3JoSlBWU50CuAVPA2iplnpGXobnjaly8t+J0U3o/JCUNL
SrKXl5z+BkmAkcqcE5gZ4GCbtEqVstyneOcFZVi6WLnLtDA1KF7SErTHHxwmfsBEGA6Yj+mriY1m
3xJdy9P3EofY7C9x8SHFJi10rJEqEyWVsU9cRs2nup3rBZTQdFDuFJknDx/bn4mK3sNKl3cGt45Q
+ArG4Soriv2eUwXGzSp7Mgr1dB3PkLDMFxtcKLd9j3EzW7plK9yPoMRKPIv67WyDGff0/bftswJw
FpzLPQtIkBIhkVwIeuF3pBANub/agVMB5/G+LuctLu2EPyiDxc9CTwy8gWT5x9PJ8C8s98wSPt5b
Vt8FtGiOZ1MdkfTyBFR6PKA8xxd/uBEESjvsKzH3dLxlUTfO3MGn7hrZcZHPfdKpQaWiEY7lLKC0
zHpWiUCwDihZGyczWkA2dM8/sFTqDAvuVeyfx6+G4iqietdnFoL/XpMyw2jZ5I8ZB25PYkgy82ys
TUc3YtyK5vGLCTK9MMsOZVLSEXVucfd/rxaqHgT+EwkLNVDDlQzX6DcA7JDyHbSx7rygH6IBEEnM
eg5BgSoAKgFacIoAPc2EWw6lBV2gGI81dlPY1yEQ4f5oVURYeULZqFpZRtQleGjgf5XcLPLPi1ig
h/Jhy0AAcJfdBbYyawHuIsGPFa+5nhMW7Sw9P183fh1ty5CPAyyVKPPzohVbmO90LkuTXHzaDOo5
1y6Y6K0psluhsWIZX7JIpG0BAB7Y3mPAlynIqXkfCiWRs72UpM7D0RTlZDV8zPsc/kVbTwc+jEB2
ehmKCIjcVYxSTYWDa/czUSFpkdepPRleH3gMGS+bbJwD23BSH3DyR9SxmJLKtOFxW+T2EiQxBdHD
Ka2nLFoRXaE+drAzcx9JLGrjP2Qxqtke/DpX/i2KOhGtSUA3ZZk3sIu4S8O5mnRnV10zi4ltVi7D
nRt8Qh8CnxQH0kwF/DLw//e8Uc8IwouNnvKRcoBLGVD9lvddKzza1HUK/ED6w+y+hwIrsHat9KGA
t99y520ltCv21Ir1TGBho94lbocA7u6X1vZOsR6HkJ1VOQMNFA1CsJRZgR8fc+JCFQTC1ng/GeIi
VjWEoVn5J2h3kJqvbqR75azdR2XheDYF02aPNGPhlBJCx4Njx4eHrxzUboubRcliCZbD97d9YjeO
2Z3vkM3YV+0IpnvhlKbu0PjLPFt0RbgircurR0za3yjMMtW6coBLhOipmbz6d5BK4L2OJEBOwHII
bOqxTx8mpTpu34MEbSUCFDiU72oaW4nhP1MFTcxNrV0Rh5Hnc3gjJXOOtL6aHD72zfXG8qc+O6DT
yYY6uKsnYdKDNW4FdoYPFzqSIMoORMKlyFghFL+RecwqpBnehTt+j8ir8DHt976dtcySUzpjfiTF
zWztZ22K1148TrJloZRYL8TYYjFsv7jzJ1u0X23cqILJZ8qA8uPpiXL6wR2owUtBtBgJ7vV0q2El
9Y38uPzC7gTFufczh0u+pzc7hCnx2dqqvEshfYC79Z5THWY9YHReBX2oVdxytJjndXE5vZbNMj24
RHrCKhPndPD/krIPw2HBcJv45Rcch8ZPiHb0yIsEX8Ah5DOLBNW/E/l7tXEmLYByGcR/MNWQSeSR
cBr/T0C9q7eTmYtA0/Diz6S0LW9QFeHYiLj8unrpQHDpPVAdpagkJp5cfkebYMil/Y1TPmJqZrhA
lBJ9XGN46URVQIY5nXpOwyK23UP4cBzHHE2cty8mlTJscMkUpocN22ehlumQmyE+KeLgZN2UyJ9/
gQL8lLGicDd47qRT7y1R4+5ec1Vppmqow/e+zQwNxMmLIjx7dx86RwPpfNXOc7Zb4ViaN2TUZeH9
xX2z4UlcmNaRpuuC0ZdL8uwkQUqyt745UdNqXFrnDptHwkR03cA1ytbs7F/kEflNqvWEP+JX2XVh
Pw3NwdQTO0YFEJtdTWtj977zlzy6XUAT5Z6AtfL869o4XWD5ZtNkORPabn7OMmQ94PNy4q0tLLy6
A/S9v5X9tXZzhTXvKLfNGW3smdavpsuxYBXbkOq7Rx2e7/hgwafocQoeBkbbPd+1YXNyWzJyVpI8
MsVZOPhkPeigjvBOZppqEFcyvGzepOtvYjwIAwLgX6Pg5eqCoo6GlwLS9vwmppYqqphYSpS3/Msj
qaMV0idoraEBytU+6/Jl4Bx2KR75iN1DMVpYhBjWQRwGmddDSBrMSwT5GLPBlZmJGW7QAWe2fIP5
J4F+2UwCkwP067CIAyPBJcDznjAA6yGxZ9b5NnIKnK4vd2BhImezB8ohAmuyb6rxrN5B86Im7BBs
O9fBBdEsuU6lmbLhJFsvANQksB8+QZLDUefcPPTc94fjFB7mQsyGHdrq6EATYFA65w/TTgbUqS/D
xwPZPnnP4yV1lZsxl4l88V/xuILZ0ErQnweqH4orhqfUepnzYKNIqW7Nc+yr8xVYhltg+2jnM/Mn
+BNepVmpYiGH5c7w4KyzGlY0mttosSa2H2L6hkJnZluQWQ5zGWSxJFO27boSnlVsE4Qa5bRe+v3N
wRm7QJ1z2gd3tyvmCkdFPqj6rTjSdbvUSWLVWUfIPSU52NQlVJedZ5d0Oy8w3vu4dIB6TAFa26Sb
lGtF7ZbCtA9MAsPNjbKH0LypmYBxNySbLe3qZZjHis5J9NVQbFhN95ytBNjSh9lxUCLI3ocpcfWx
XELuyV2QllOJDQ9Om+yKJa9GsHFcKz1SAUyxcOqfFKbn1HXQ5l+Zpz/bQ17+7bDNm5nQx6RBB+np
935SKrBP/zNi0AEHYomiStvloxGmSs0IRM6XejJkZuhflxniyJtmH/t9fX7F+Oe5R6jCidweCUg0
JtFDzfx9tZV8OXu8ZMgwtOpvBsxCivbeJimRGXZCP6xJ1WefOQIDyTGbDEARdNf4AUSNhrFIslzA
rY86UjTPYKe/ZWDsxsSLyripPuLEbGj0I3Tt2wUQ618fkYXbn18JfTKY5k1s5Nmg0MZyuVTccL92
l4cCV7V/127w4LL1CNcgVhYmkDBHcJgRw8oY3qae/0JA66TCiT+SFXJPNiCE1NxAYIu2CFbTm4yd
9uFBL5ncXvS1Np8fnsg0tQOe3L1SADauPQypz8Qti6B4s/JM98maPZAb3yGCwnJdC0Z3xaCUq0Vh
KtiOKv8K2K9MPRXUZwWFmbHzoMOvLuvCZ3U/Bv46DkCBb0Fik82olV/0lDIvBmGtpIFwPjQWOk8n
Z11VFotggYBYznqTxdQUmqivsE1sDeld9Y9LXaP/KTYEAfZGnCxQnXbKgPEAOT6Ispp0vjv7kbz5
cDVLtAjTNNKr/RNV7RERvA2i/y3X0znX/RMAf9CdLhtNVtU0LqRRGmmQfFL7lL2nkcERMUSWBiNn
WVZWmbltEIArJ4DkE4VStj2tgtHQt8ILKK2dYIbXHJLi9LYVFwdy9VrPquBFiqkM6tByzmeXeviC
MfTtHDuZJObUwRC5rJvOfj2xocX579bRljLMpn/IJor4dYRI/QxuKGAEipxZbopp2wZFLjAlyAdD
ODtLcREVd/gcQTH93+tS//z8Eb3FeeEuU39/uy3zVQTyiuBp+CPBJuBTth2SMu5gPh0B94TWVLok
IH7VrFbJKp46toItuuBrRWnXgHzUHFM/Jiy0HP8f+XsmXyONZQsLeFW70uVKrK+jj083K5Q6SWej
nASZeOCwfiiFrAKbzUe4BzKqexOiYsJqZRg1rAYDEpp4OgxDVBWNbwKj6XXUL96X834XrASHv0BE
y/6VxeFsnj3ijxJdpdI/YtAHCsX6Bgk3SkNm2EcBrI9GeiXBHt0oGaADhGf8VjiziY1e3hgItT8Z
vY/cNMdwkotD1nqK+xFsec8agwj8Uop0OuQDSvmwveNdaWsDfSAIsYkFI+0DWh6LghbkPQQEVv2+
qjbSshq2ai1RpPNzXTUCM9tmQRIVfZGjKHwyHteSXDg+0TYWVGv0+LH/qcsW9d5ILT6cdGYi6MYD
mU8uZGdPSSy13bX8cvE4LX46GVptpR3De9XvW5FRsHfIw4+v+oniOJtxoj6uNjww0bnoPbcC0R/R
gxrk7TeNCORAwU6BIuID9tVdfjARlCiBk/Vo664fZ+UeoSJLX6725iTNf6XTXIcmlp+7VEj3tC5c
ChhO0wNDv6q2VUXtIEHptGpqhDEIzrHKy/5Kyh5R9a28nysr6Xoxu+9Ax/4XNKbAF/PxOnHKfB8F
N9zRyVOZAKaUxEI1tMJgvt+1kubeAQyiT00J1i2euSnbQdZl8dgtx/S/F++O29LNMVo4/sIu6OIt
ZySXynU8tNVxI6vXYdIfeDG9NvqxkcoD8Pr5eTiEJETHcBn3UW91sSVoqGp9ogFch9IqTatXAbCG
SiooTiPUu/VmBQ2ZWDYnYDOzdAqA0zkzbaE1dF7zyqwqTBI6LzoHlAGM/LL74duqUn3SgUJxb1X8
tF4+2FmezmFd8pH+XVG3SkiG0bh+mA9dWnKXDoo6H7QhWsnLJSapnL5Wel5XOeYz1mIDQxAtecm8
INRjXIHjIQV3zK9505Pu58Bt1Z8sRGkJF4iKHN5QxqHROSueQGoYuB2b/uxt8Br9zbRaJyEU29mJ
VuMHkimgt0g3MABJ7+VdmVf9n3R9tkK215XJPW/1ZxX1ukRJxT77IIo4cLCbgBle6TZfyzRftNtm
5RenrSNw29T7aFny9+GeeHNf0sz4iEy5QR3zvmGTr70q52Lfn+iV8MLZRsogEs2PXb1bL29sFB4t
Kih5OW+PE2aWAI1WE5mqe++jcW5aJ+Gs/2afGaCZYMtnYXtGD7UJbR+dSbQ3hmQFeXYIl4loReRp
Lu2fqa2gvIJ1FgDzcmImnIWOBoX1NtiJm8LIdE1hc8pkcN2Wnz6beO0iaSIfNBvZVvyymZfVPcSF
oHf46PGw0SA5QzqzhItT9kq9zXYSh4RUyMHT2IHIrblcBDq5SBy/Ms62mKSZnCN5qj9tNefyEczo
qL3nopD5OGDCd20hWswDYvD54vSQpnIn+Pl5Wt6kbofh2idvfY2hRo5/G+xZZnKzf9QGldb8aXpD
loGOAM+Ylct1mmMxcVNCko7e8uwz2rU7g3T5aoq4CeFLfrv/mHrsFeTquWe5CLnceuXVnf/rFoYu
wDQrJVo2Oc9wxszIRaLtTlKwq8N7HF9hmiUZY3UrFRF96h5gURMPwyqeirZ17Mxp4KQrKSl3k+cw
8Nd0JbE6t+ZI+EzDqP+aeW9GhsYROLNRZ7RpSFTgnw3kQ7JWIugm+4X+MwKxlQY8K7Rt7LJBoykP
ydC54GSvutmFKkHIeWfnXG3t8VXaK4+8RysdWIn1i1BkL7SPCbO9yfRGPsm2HiE8BkOLhELQeUYz
n+wiaOVg+75wBYbPOuH2EvVneloukfSTSu5I3mxHHUZ3r8dagPtALfR9CS8lbnv9wbkhAHHG9Eoo
B4M1BEFGhxYoKLklp7oaYlk2Z6IvuDBWyQMaG3Y1gVPnPOUD91HV5xenrZDKS6+U3olbTuhoNy3R
4Rcyx0D2Yllg4aJACgoHV7OZ7g7p8GOUhz4/6EDX+q6+xrfIaQknt9zdjVpoziyCqWVp4XDuIGJs
os4rXxdk7Jgqujz5OXSVvt2Ur6buqzOZ1vyEahbyd3u2sMgv8WpsCwBP5jt8SDLiTPQxQk6LDj5t
ni6h346adHuydNWhQOhWojd4v2m5mNbwGI1Lxa08ckxM3tRfQB2wiI/3ulIhYzcZaGj/9WalhTeD
GfBrcypgNzts0yOxJOHMX5MJP/LvNbwSt5G0fvsP8zwS8opZj4PuGAm7C2NmE9w481yxZnX+s9oz
MDNMMJEBe4V9LEq7+aREH8hwty5PG78yzpTZneth2rUKm9fYzc2p8og+2kW9DwH4MLH9P+WVav4e
MjbtW1D4bLOIt95TqS+2M6kGVEW0ejauGno3t5ZdvBEKm/aj599Bkj3zpIuUcOKkPepFmx6Mcp0C
NQbgakVh6Pqu05pw9Ko8fStHwqIKg0aatIcTNsgjVSQC5wfACXrlNPro+ADo8N1tfiiIFAUy3e8e
5hHGnwLLhOjtaLrsOqDOn4nXoFf9tlfC4jW8ygYoOZgBSPsl9gqX0IOHOzWKhr+BpJmsLcjQF27P
28HeMwsibqLXHJBoDRg5bFOs6/Nk0gKwnk712X8DduU5NaYSeMrnElahMq3G21Bu7tRaLtxzPHAo
7bR1v5bomhG9G/+5tlAJC77vASsgex0lQ7wPKODOm03CeYtdvR+l8ODi242e1V1MVBCvrSiff+X2
YAiYY6S6MfPCvuDPQJL1xqT4AW28RfAL1gWuGPOFNB4BoylSBxvN868DkzA4KItlIFbYtPIe1W31
EOVu0P0wu344NhwDkacoGHBUnVfJ1xzW9eaeWSF8qE4WXHOl8fBy7O8nim1/H+yEsndfIC8F7nNy
ht31IbqZvxznC55aEfJONyMgmUkJNKykn9MHBfv9Ybb3a9ql4OvbQccNdlVbfF74hnjViNiZB8ls
amr6d6fXa5lhmWeBIVO9KaN2oHo48Jwq5VChZX9Me/xRr25moLdHBK1EqOgiraHqBU23xoucNwwt
SoLG2P3DIJF7U+ubpt/Bg+2nfUBp3aeMOZ2IAEUIYKQNfoW6Zxiujwj2N9TiST43mcjU6hnwHoso
SdJKC0OVZrGkcN7f1ou/IXxGw92+kkmMEG91orRjCVh96cAMygdYc1hPLNgCKpDPrNWrkJ2Gn5E3
bfSN6TfeQsLM7bkP/jKpZel0ijrM8K3b9d8j6H94Tm+TGi/Sd2MxgU3QOmwG1B6XGYqq8dJ1py+X
fE6kklCuN7zdF4S4GxLK2Td0SIbzHcL6RL+8MBFuexb2jZGi/UU11G9FAJ+OIinEUT+h2ZYbnWXe
Fdn7yVo4HeAVudKtebP93TJ50AixgPa98mbf/BZUR5FVb43ctmAE+tJqsS9Y74sjeBUr1IgGL8mB
bSxJgiZep5x3rDfl64necYmlBzwt5626ocuryhEwYZfeCAPnt4B2ttCAlAOM6Mqu3qspA3JRkZ7A
0H3lDa73oztCxgmiiGjMjPMbzZAQLCBCUcBmBoHqWpkFPUrqO/ho93qSPw+DCmwxbB9sqt5siTkN
FUqs+bImCFEg64op7ZvrCuSlqspT5wX0jtMC0oirqvUNQPB97QG0kmbUmhAXOFSNcnwHiGvb2+Wl
PxgWLOipDx0p8/e2dcQKo+AmhbyPkFObxptPTNgtwL9hntu9GzNane1/7a1KuRNiciyArKiGqevc
SDo9rC2H1+QJQuSX5PJm+8kkfsrMkf8xaq8rPDjtx4Yysq7xlSMLmKLpLuedh8ks8wuX5vXV596f
LJ+yHD8pkikstJEUg/JBBxX5430AbnAqI4lXNGlBQRnMbrtyW174gnR4jd/hgmCE5bXprsoh3lZE
1/V8sg6gduhY6fWLjaHq0uo5BVvrjYlalAbz7I5ZGinsffqi2RbO7M0zWz5HXL0fZErZKfyQXBLF
bMpobAsrZLXpzmvikgkhhhKYlKsbvr+dXeqschDq3mJ2BxWnRQ7fe2v2VIHBWTddv2zdUavdCNgJ
ab5Bn1IPOnit9tW5piB95NNtQQcYFG6UZdtc0s7rF/9DUe05Ahq3pcdyjk/II6NIZRjNQOZdqDF/
juu+yorVzc0oKf70Kw1r2oxULSHzHjpN/VTSQUpTG2DXocJJ4CftdJ2sXl0jwqCa5HwWmbOsmMwa
MlBZLnB5TmPwS0uu5bv5KxXEV5YUhKyhEaHbXkO2e4sXTcGniZEA4SDF0OHFzwHEG10WcSwe+Rla
vH7MT9540E3bjgZ8VIWvi1f5oLl33VOnvmde8BwApTyzykAhQNc0rD7raEL+p//zmDzBIlWLF0OF
N2S6MyNjSUdJjHKrCTyjFOY/zhdTYoTttDpld/ZCj+ti9GaCKKOEOjciii/NA6avDl+kBU49pn9E
Sb2AoOXo5ScnRpESGFp0LnoLTwQETiYt7Xl7OC/jq/bVUWJOcNbcTBIHEOoCineHaq6iKYdza5On
+yQZKBxQ6quQu5F/Es/enzvzXPLbVPrb7Hm1XwuPQ4VJZn5RruT6Z++eT5+43g+TlCtWEBBYfCBz
P4Elu3VE45p/78qh+RV1roKctlcvDw7y9RbOBcfIe6KD02VO10L1KnTzWJasbLLevejX8WyHnKXC
AzHZIkOplYNrP1j+3wVqcKbwIsJclGamxxj6oyTV2u84S1ry6Ek6aGstMihzdFc9zEsgpAaaRe2T
IHsPOBVcVtW0M0b+t9Ov/zcALnDeu9hjIFMLrwLpBKfRqEz+Lt+HbeFL/GaY2IVrwgs8uwtfxq06
weC6RsVWiCzE6f0/hcF6sYYTC2cAE0LFbaqtIa5alwMdKXMAOlhZ705w0IcW2a1uujLyFZPLcAup
P9VJxftFku4qNrC83TuM/GCCO2fZt6I/hqfmOZ3Ob7SpY8Q0ko7gEMywETY7DQtd5vle74SHqAnS
ydnJCVLKjIb+ommCDoZdNeUCLkbREZUWmKSjmU7reHNm6SznxsQdbCjnjBikppF6ZFxw+woVF//G
85e/WCTX+zhMRn4Nppa+kw73AHe1HTn9eKVwCLoshbRPiEBV/D4w5dbIzSF3cRkAjf5eOVMYCQFk
LsRcyfQDqAWc/ershHreqWjGq3ssAN8h/RtLjPrHR0QHXaehaF/1CB2OE4zyEuSURqiCS7k1ZBeK
6LOam05e6z8Hku92eEH4UZwyKUF7c70ZFqtnsai3shxeTauM+vtdKQZ/yhDk6dL9Q1pO/RUknbOj
vbCHsPJ3WtwXw/og2WNX0WBhAZ82/Wvg4n1gCKxR4qmwpUo0JrIIvapKwR+tC5mCP+TTlcR0B8wS
+hPb2UcmHmn1bM775wxqbE+kdr6xjU6Ri5lwwxa3+m6+to1jUUqP2FCWeTCRqzZ/015e7JIQyWnN
gcoADiYNl17BJeWEUvXvZICv+vsleE4E1ulskkmqalztOpt3y1/niOEBQ9r7A4ZX6V7VSbs43z4/
Sq8y4gIyJYo2wEjV8Ngj34+o5QJv2NCEtnmzFBsJeLfjcOH8L9UHoF70rZma8Wb9VEI6IRtMEc3v
scyjifASCXPp7vKKa0ko0Y9jagvroKP8YSyT5CWVAof7kXoQicywJeWtA0H1eSVttNSYYsfpiP3J
fMp1m4zPB9uc/WPv42BcxhCprDQ0UbTlZcFD1IF8HyxhI1jUcI87xqY6dQjhEEfdwm7VC/OhMjDs
xt5HM6xNTPwiRUm1sHmVp3Ay5siqY7X2W4u3keoJxca4Ub3KhedD3m/E0MuF4NL4ZPcnpxTddH/X
rhFzc5609ufsVpIZzZDY0B1kzzuOBHmV5r2KZiDeFrS5E+HvK3QZNFwc1h0/9O70V9QFhFo7Gu1f
EbayMKBuKkODQ6LytX0xM3+6QXTzKUgl7svzUfeRGVj+JmsHjbQeEqY7Ird2TjPq5jTP8pnGNicX
OC4IXMFBVr54EViS7fzLfITCBDN5lji5zFMtGLKG2GLVqfvLWDqlnCqq3g0b6GT29JZnTOiIPeUt
L7mdRRU9ljbtRIJgoAgRF5KRxLOzvZfaeFdki0vPnY/IoaqFBpC/7DBIUpgahqp8CFqNSUyTbaRO
38xBszRJ3Lb86FPJjL2pG5H8eUWsU0l00Y+An3sskIMVXkjUYgVs06ZWnGFWyM+8wSPNeyCAHtDC
31iBEHUUen2FD+qju0l4tXBbRC1yqajTwbFomP/xe/1UYhZCvC9yjG9bBJa8xKIjXvavqnqlkhz3
HsT6Cg58hxs14onbpBdkM6izwx0jcESuWxi/GPAI0uSok0V88GSDWmkUgAFP5qJN1nBrSZN1HcIO
r6IopVzSjdi7EXGGOx9OgYjLDDk0q/RUW8ABRYiFnBBmTEAxhv8HpYXXXp+ywSY81Tj5MP6f1NQw
hH3Bae4hToGiMctpKyH/NDIQQc3myvXRWiGGEkEQt1nsNf4i+uy1+9Cb5WZnN81nkd2O2FidCQeF
JaWPUuCfvCOk7FaZUTPT68wJ/6by6Q/zPQydfKtK+UalPDSGXMLrHfRoS2P0qCwFAWJPyL+mMtQl
4yLx0/zECwV0ZDpnwmac1hUqWYFyaS6tbPrth5NiaBccKlW8UyZnbvw7sxu+8IIhxPf7k7vSKlt+
NnhXodrwyxsO/ibzFR6Pe68tNtQH/j4quCKgoUPdSF6ZhS4uGffaQ2vGEWR4p10wd9TkeyBpFv0Y
5NvFSwEhIMRun3meYTbGTQUIBosbBrEgbCCSC3ifPbOeqRXK/ozxrannVCDdYRbl4XSnIL/IIHLU
Uhp3AiGvCvTLBQOfM1d+KdPzlPtg5NttYMRqX9gx7/KvVX1myOkF6VP3yc58vbLK7rG0B0pOO55v
4J99tKwkp4wzUerie88uBVmIuA6NyL+KlMlfJOzcbXAqDGWrFwF+nuLUbgXpJTqnHB0q9dZhCHWI
rzTMsrBaisRzLzPEZfT7szm+NmYeux5PMwGbzanhFf2ZpdYLUM9GO/whHkhk/79gibSe6GNEEZWz
QBl0SVnIb9B6TB44iCk2kkj53xgl7nINcFGdYw9K6wETbx7wWI/8bdXsK3XllcSqCBaSLJWjSwLX
qUB/XDejLc/QAQun1aqNCiClfzyxkZ/RpoHZ3ZwqVLt17UBywj0+62SllsrqGBfhPdrP6wgrBR8n
3ha79qz2/4jLo1RJaFQHVgDEDFEFHabUZBI2R16IRRlFh53AHuPlNdc1mxxFUYGItwzt1WI7QPJ8
aYQoF1UzIa6o+VngiOfXlV+IqDlMn2RILjvc3MWBJYTUOZK2URQvgFdJlTBjuAT08nDb1yqKzus5
lAYz9IA0oINClPN0I02Ob1Z2X6+RZc3WSitV68qq3qKhqYCxhiytpPD0VMlzFVcqTlTstWTyl/d+
S5b3ZFlP9YfP4hbXRT6Q7m3rEjTeVcVY3H2xvNVYXZlPngmr1b1mkTX/oFB5W/UBy5VpLCJJ8puo
i+V8b+BmcZmADlr2UniYRY51t+Rm9x/q23PoyZcwYbDuEEbLQLWX7cyOgoHXCzmHYK3e1SDHvKPr
rjgEHVsCWx6jUJXQgdCtFpHRziPpZsah1fSR5/8xG5utVSwD3Bzxf+QnvjouihH7PDeNtG9iWBUL
1Wj1NhpS0KbqqgIvfc2yszxIAPtI2Eh+wMbV/0/pdZPvmhmGC0yIO5LHpJ6zkrBqoTnFN5x7KWt0
gR6QUGQwANS6n495lBs4cJHqAjhcAeJG++TmctlTabG91plrK43J2QTnfF0PpUXaDGWzWSBm3RsP
C1PgyIhN+yiezzOmYCU4RK+3AZ7HaDJdvS34FfmRLmpVJi8fhbgz5xEOvN6yUMCzCzSDDFc3/g0j
/TjwNN3jalQMv/JpphNWrlR/ezoD+MqNNTQA30PNuz0DJhP9/RLfOD9hCybsqEIDZXZZ0XNUPtgS
YXNhkmiAdTlnOEHK5EOk6VzphRVCK6utDRm5zhhu4IWY2GaAniG0wXnFRG1oA5sVVD+TJnwPWGB2
N2PO/k9HbP3Q/3QTMFwvqa1moKlodolZwYlypTmJBen17GTJ3qihWsJymamXPAaVwevQ1VkoqpjY
nzAFjVjeGrn9x2vHFckJz67uMhxiPWRlBLI6MgHSQpH8PRjosFhjydb+Io1YvHMrKxp1bH4vSjNH
+TYoZUork9nupPKeDpXf2K1qImvkUbvF1GEM5OnL9h74DQC73u9G78zAZnORqSvmJ+Kbftld2h/K
WaeinKUwQAUVAZ3WDU4m0Rus2O4tDq/lzqCyt9D1lPxSz1PAGUHwCnWz6O82BuozEeNmWSn3N1V3
uh3Izmpa3DZf6WR3FiS8LwAyrKKHHd4Qf1FZ4qy2AkERZk7q01XF0B9Hk/wevMXuFdDOAiCDz5On
EUCWwGqcMXFLmBG2yIT3psJS4i97SAJylPBxFQxnSk9WyEP8B9DGv48brdNYCL5ei5aTeHmeAdtb
u+sb+EDuG6q5mk8L7RM4xOjkL4kjp32Ife7xkLRX21JGib+LyF4SWFESTAUJkgV3jNMCJQggP7Fc
lHosDzt3RvP7Gt/3OztHfhMvzvMgAO7vdVZ6BE205avs63gn6leL3puiRrDf860/9g9WguMtQeEP
7MVLH9BtcyGPP2Wf9rJPqcj3tJfTJ8uko8iRAN0DnpU8qkO4xgnyAiHuj3E8dJ54shhDe8LRU/OG
+PRfS59X541IEHu9npmbpo5n/IjFu3+ZvIrk9KwdUflAHj9Z6H+wWe1XFZ8zCXsA6/9lZWGb7cLT
djNTSpid8IKCkqasmcLRAv6o/PAl8y0sKmeQIqfg+yC5Gd7G80f3yJ82so9kQ83lWEaogs0FVQMb
hjS6VpiykMKhEcXmJn6j49XLQD5uKIeIXjTSJgQ+PQ5MaLR4cHsunGf2sTzdoYHG5jlmjmZEBse+
3JONAP0+VZQRLv+qo6XZxGBwzyNsqWacKi53H77PpM7Tq05K/tKuaCw04OFQMI8RBUd67mPA/MCf
pdSpRt1GINpuafO+YbzpU2OhYsuXv56E4czuEN1+YDTjVPqOwed1dckxDl9bFd9Zb/3RhYfOIiT+
6E4m1KAk94UCSwe7FCFrKUvGi6fxlezWSVoNsne2aqgnTnef4KhHKTupUjLewnbhLGAdhglNAFRJ
uoHhrn6qOcgDzaIHGKC5a76B4FCWKPripa8evf16uy89RrwuifkSKexQQ+Q6G3vu1QcLh4ziHag4
yxaDdZCqlgLBH+LMnO8gWTk7YYNvwGkZQrzXpzF+7uwG+SaL2xqXBGSVdIhTZUhPDQRRr4Bn5SrG
7CE8z2VxFsFA41aWRlkKFrpkpFeUJL3QcJXqVn4GNN3/pHRYnLcFuwyNXQcUSI/SDGKbXoytjTI1
GToCi03U0BlHA3zDezOPQfh/Z8Zlb5BIlV+4au8LWum1sl20qbK4jCTwQGXbV3xv8IF1zPlWsMMI
2a/gqFenuCXht9sL7ZzHeL7410HBfsDdE5+glar7snRcvoT72Ud/EbBePe4Uh87Gpxti+8/1P+Cf
Mp36u8qzCjTF45OWEyJcUyshMHpx1GkBty0nNvlaElu+E0sYZuAKbBpHp592dyqn3gJ9PnnVBBdn
W7qsmgH/55qJLH67/59TnGmd2dXyBGZZUuRdvuxk6HbXWxQZ5axCpRlu2OrUGTdVeGNLpRgBai0b
xqQGMDyP3cut0TMmOrCTOOhLbJN2g8t29tKKju1qVbcaNSGGwraYUunKAmJ5sUeNeyoa2HFOl22Z
tEY9/6+j+Z+WlsmaSF+ayVEiwtAK37XkNonlRvhN31vgOaMWRApGPEw6P/OxvH0GpVUfLUWdiQCI
Rd6d3dppcVNKUqstE4hWKl74p00knseiDI+X66w6ui/sYKaADp4aNLZyj3aPcX9LeAkZTk2BVem2
wnc/Sb2qNZUG9esazgrE4bGdzPd86A0VkxSwPBHaV16i6YpLDcHz88OsC9XGNcavJvZSIk5JjPtN
cuM7ftcixUGf+4mVf+nkqcXvAZJBVmUbSTmeLDlHzkc39HjJLKembyfdEwPpzV1jqccUJQm933NF
f/ETXq7Dw4Q1x6VMqUgbuyoNjES1tm4XDD4nlmQ1AebD7kt3Ym0zeYwZrQDqe01LZ9TM5VWwjDOg
d41tHigURqNGnVHwgQPstwoftmOSqZnNrGU2wFxtH9+y+0MGsV9ySfnxgj3Mx+XDxv8zSlByfdnK
fYfXNW2X09dV+FnDU2N3t5FdXM6JmVZW7Ik2oB96jzSp35Eryimkg4Di/xXS0CwUwdPzCa+DaseR
2IXpEhq6vqC75NmEGiuO3lwncFG5KrBu1/BQM7LOKjsN8yiX2w78bCv0Zk9mb34ULJz+puV8jBEy
cIov0XVRFnbWihwrEwUrcX/Yb+F8x1+iq2z/3uCDw2gslclWe9KcvQU2GugGyV5tZLVQbpBz7NbR
U9fpW6vQFaunl+Ikc++7FuE7AYAKCcbKsbe5i3/yJPKsI3546EjaVWrhA9QIFcVvCIhn9PoMmB2e
8GKHtkYq1Pln1NBU4kg6czQaLq/UZMqorEe7Aw6Xq3D1M0PTCSqqVdyFZ6/gmWBIKSwIuQXl/4H2
m510yWDyyAy+dm1+xnoMMHuNpvIp7WJ+ubq88OdwTwB2mw9Voakap1zdwUF2RHQqFW8kZS3xcJuq
rxrvWYho9ez8GpJ500vYILGW0VBGMI0DgsGwBRfU5tHNP6WtesjYxoTy9657HMY5Ia0SgZ7UnD4i
0NsUwZ1Yo+I3JFDFijM/HGzNpeArzploV030sh3i5jnC+JRdL8aIpxnBFnBkwrAK3Wohvy4nQIpQ
ckaONRrqj+TGGIViw+1JzzGAc1uTZ4cnUcyamUcVVaNvdZXBK1zD9H292EqilxcG7qzT94udcpJv
oYTHyKCtX4EmUQDdYLlSzo365pyonYhorfRubYJThCQ15ad2UUofG0Lyr+DCOAFC76Hg52LG6qUU
F5819qhgnDlOWUbk7q0+DkNqMyNaGmou+sVLBrs8MUuu3PoTS8NYCOF1Q49gqy9WTakFFQasREQ5
mGegbm843x3xSk1BhR5j6K1h7Zr9Kv270jopWv2FTa9Wan075A8cIF/4X1FLGWEZ1s1a8xtbcdsA
P0FrB7oFLvGvCEfMuP1I0I5Z9YgPPbflXBo4UQRiRPpWHqjkGkjF18dPpVksNuZfpqBOBTg8xsv4
YHgpET5UCSuPMp0VR8OyPBroUWhgRUmEK245Dxd0HlP4frmxQESny6pVqF4sQ7eS+kJe5m81oiiV
APYjXFLstgEFFgpzbmQe4po9IlaAe369phTpn/8GE3s4awrt2BJLFw8CBK718BSQkUaYKwEamCMZ
NcdQYqKSyTJBu0W7oUXSYW4CI7qv5MoyCATLHadcJMHIyBtVF7LuHHGqIdc+LmN6N/CUqAkMD6/V
vlZCE6VmTChhEY29A8GHotA8CrAPDhzTbT1fTQAR5fAxaLzk8SEeCeCOFVHzzuZH/YmCqro7YPB7
gnTvOchTyqB4wjYwlje805LNU4yDtEQMyIeP0Fq9oDjfiL/OkWJZPdW6noWNZML8aOLqzyI68K7k
UAF5t/HOoJgu++RTHeuOUxy6RTNCtcaH6oqsp/wObal4OWgc7F+NzYIeowPdUtA3oS9AwUfTXsO/
npawQB2OLfyJCNTKhXE/Hfg5sU58CzQSSqIlH2x/Hmy4Cly9as2Ckcb0hwk/16YMDpMxqHgN/30C
WNMjVMy3iApGakh9s/v2/EOnTdpTFnUH5Obymm2OYdLCgiayvcHuOAYdoDlMofUN9YElW10hY1A5
0gJ3MK+nrsgvIu2bQ4pKLpoErOz9i/H4p2GNFuUDM+/7sv99At+uYNg3NaHTKv3CDIamDzcPS3wX
prPk4mHDmZSBJ4GV3lKdtU8d08Uz4LwtzyhcafLCii8TjR5rdgDTGg5DyFNZ9AM4fNZgIpKrkGWF
8O0QkIFiyU4jNcSQVp0wLjcKkdbpiCHXGvBRqDVzCHXd5I/XLzDeHwe834PZjQSomRkj6ulRY341
HZEziJNp838xqtsd8IJufExaMg/A+Fc8AwWrOyQ8MPjcRcTn9UJ0wjnCEbawsY9vHNMmJazrPajT
wj9IY+Mpk45VJf4fltJeEt5k7iLzUeBlzmhXMYRmESOMtnFy/CAjHfvUXDvJZfGM9IZ5/TdbX354
fZNwqAyS+MfjdbYArURqXQ9J2V+FPOW71R3z+dDtLId1XKKflGGyAzxfP/GxsNePhNHW+vMgLqQu
N0hdSO8lncHmRJMQoq6bzCs6orB5zG7DrA4q0VObfRdQEcGosepq/8Xhy9l1wgmZyoeIeWjTJv4w
94bAuBsa/t3krPx8WLN8ZLltZ4c8MrcwTdVbPBM3dVMdO95uMtFUyxQQrFVsIDJC9PmubiqQrU2E
bDH52UIzmaySx4b5Hgu2fhFFmd2HcFKCr7DnhOQqNb7KXME0U9Y2/qfDZw/u4VEpMHEwjyaZCYqS
AB4vOwoEpeCQw63gFEPyohoXN2VXFGQIaE5Fip7yUAZOTZQYftrSrbYZqxhQ1dIvNuhQwr6/RmRP
MuP1aHu/BAiy2RWf7Ij730fB9m7m+fukx4vD7uU52B+aMyU4X9A6DSg6JUQBeRm75b71gnVwSAGk
hGm5GiJZKmJf8GoI2VJ4h64GGhdXVTTN/b33jjV0YgttGkw6i2Yk/bU5Pqo3ku9vBLua39StQtEy
jXGvBfwyhrDxMGUfZBrkpAgJW0Q3SX+6FdgA0qyEZ2LJCrHo0CkUAIOtY/0J8PtfQFYtSKO2Tg02
O7t7Fv03vwl6FXJQzecWm/uQyMxFnSVcOaxhP5oI5FYHBk/bdXoAoCZBddEfLgPd8EnvMZUlIEoZ
c9koGAZrE5XY1nQCD4zTGBVg5ATGUk5nqwNvKJ7GOOkCIUbwhNt5stKoR/9Z6NC/6PfYpzkzmyf0
+pwvD4ueMZ1s3wPf4V+VVAyeZ96HLiM2AxSQo3bsiT7otDL9R15kIQvvAenoFxT5oHBx83Jf3Rb8
Q30sJljZYdyT41kOJ4Ab4TU/oQObQV9pAqlLZQwYKTIC97DCApfAfKIur4NDq1jBPn0NuRNPQvOB
UFrgrjqdOCiCCLiIllgij7v4xFBDVHMDhS+I7xdjNgzhcuVJHaufUS1VVkQA2re0D/mNUWeOfSOS
BFAStlRyCrS9NvfJ63hst61YODCBgItVo1VC9W8A5hjleDnqVaEwJ1YpYrXftQq3fk1ncuv0yp7b
cGgR/HIAD2JmSCdrSwtjmVwBO8IDEGt+BtBMfH0RsEo61BkVLroz/d2OMGmrGPyqbkqpnmPcWVez
62UyMcudr6GrKmMG12QYGUZ2PzgLy1/LiRy3aydGMbQ8UFhw53EWbHnhicdLm6wqIkY6u+uAlkIX
WAogHdiiWYxqd85zlukkAWv/5O+YAy/7DPyx5moTo5DtdLpe/r8SffLTyTtE4fWMokw9Hwu+mzOg
iSYrxPBWWJpW8pzZsRc2Dq08h3CeHAEdFRKRX1fhWNuSNkvci6K1mp/0le3QWwIi7S9gzMJLqDJ6
GPACJ73ljja+0vSfzRhoNvVTC4ZoS+KXRkWQVXXjwhEgyMvg2egBkNXotQeIRu2Dy3rnSxpSVRou
ATWclLprauxMpgXdqv9PE3ALgTif3ilxADT2X+iG2lGeQW+2WKAdovsfmHxKXj70pRD1DpROWyzq
FJG3JMYiVtToxapA3nlekxve5LKW5R9sDUJqtEslmqt2ZyzdSlBUKnirjIWC+gSL6SZPeXsnNxJR
an3fueteo9VWocfliKQ4+ShnUvw9P79U5h+1VBstWGHLbkQoP47HKd9nPmAjyXajlpru/GEHaO2K
xe4z08OKPaw9RiAeC8OZuQBY7z8CTVND+u6PZByhwXay25TEJe/cJQD0Isy6EVbwh7x75WB1FFeJ
w6I0qn0a2kn309/n1W7VqwIqSSF6NPNFLTISYTAvW+dL6Q2K28EC+zSlRqffJMjm8mf6VCalntJg
hsmP86SzxEq4LfXfOzRcyJFyj4cPlSKtBGJJeAyTfacQP+UAlvmVQB2yYtWDHNEHzuuJqySl/MQO
v4G3z6F5xLq81AwcDDY3MuhLdBYWxXUlfEqxUa5JCRrf5jhGb2Ox/jukyoh79ju9qdRqlyltR2iw
3A1a3UHgHjoDRvyHADaNWkSfO9lM+eu0C5/fDmgFmrFo4M9d39nej+bKuE++/uN78hFtRf46FSV/
E0xcF8o980zSk5b09TtR17Fp7B66m5PW4LRNtUcdQw8uc1d+nzuT3DIlI6yWunz0ocKTOhgDY8fK
sjwvRr3iF/XwB+bwQ4EOuc90bA90FybbgfJEm3qr99NiWx1QjwwGFqVfiUqmY3MnOG4OKeRlRTHo
XFce5F+2EaP3bOwEul6adWFwapXE2sXNYEe6mZpPivgPYsAlb5nBdUAhAKt0Vx9L0mIFbFGW0euT
vtJPnm9rH3xW4AbhkmeBqraLEo5DZOb8sEfMXd6TpRZxTtsnS+PtvTXWNL3cVjxXmOxO7jyZsOc1
uK8+FiOAGqur5Nm4UVN9oQCZqN9uv2q5dkjYjSDFcYMTSF/4AI1HWJY8a3RjDtYNZQb8jJhFu+Ob
SZa1KhSnIaITZo8jStiRbB96NTNWhlMcEo3nsCVamchIWpUm1KFtX3sWjkGSbNno5GNqN6KfW//5
lI8xbX9aeZxZNEGnmaxGcwyETEwcN3DymWpqf0Vq232o+HYcoYab1UnkBt7HtbXKWlHrnHs/rYlv
Eeuwjp+XD6zggxkM7/WAYqtT3ilYMggj0udlsRovbLmFg4B7Uqs3x6u+C6+Rdkbiqeub8lBbZu/J
otcV1VI8oYOPWqRVVJ6IDK3xa2oKd8EALRs0HiCjQdskqDEjrZj5P4iVFReZHYC1lV+oQO9REdcJ
Mtx8UfyH4vsB2o8l18kFQ5kHGTaheQPlw+Av15sNpaeiZC74yZYPAxfAUSRt5b/hg4M7cGrqc9WH
NDot1DgSp5byrxYCVOJxq86HovgtmYLZYbwiaX5Mi9KYH4Qr/yFcPejbzPb0ZZJKmi6QjX3+o+mM
nSJMsQVmZcjx05MS+4NkE37HmQrjfyu9I1WqnTFWGbx9Zzlp2zAYPqVPB07SCzu5gY5f939enZd9
qbLzjQ6y9q73E+my6YiXVuBSeMg5r8TuKS6SXTtGCdoj07UZwjzEnFCqdJrAp9Pe7cQqV/FPNENs
BEHwvvAzixq9GFF203GGQmY5Ii2G3XOYF8hoevP/OIVMEF0w65sZuIZ+KXX9jZ0P63aH8sVGH/NI
Bkh6rYy8PErBX3NKbYPlGZqUSF2bSAFRqgMxJHkqs+/aG5szhoguFQ0xMmfNQ7eiH12VHZg4cP4F
J4zaPPLFiuGQ7Vm0mPHMMyaMisHBNRh3dXYmdNQ3lzBBeSSso2LosPbHttpcwLvQeDEFWBJvctN7
/gDHpdHwW6nYc8XtvFca7bdQSnVn2Yyu+Rw+pWh+tuqbPSwT20lTVIxuq0s0tDFul10z6Yh6ilMK
P+jMrec9T0RiWTWAXvqAuKmKEZKUbvwoFajKECXRQvR5DCrpZFyzkS7EEYIUVrajB0q2wpldof6n
Ulq5g54Kn9uii0Wz1gxI/dMpiLlfZG5QXaMHEOwzHskgmcsO3UHihK99yGtyOPxQBBYtb2/LWnHi
e0J4P+R1z2q+2ZN90hyPxnHiiUM6RcgD2Cm1cyMb2HtRiWgTyXs+UXhDoGNDU9sBqw3C1ZIj8bSw
ObmRUniIIrKENxO9a6K4Jx6oO/z2GNX0vWPDVNVqhf2KH/IJPeJEIpI/tf6kp8WqmAOfjfUOkpKA
RwufRb3RXgKz8j3jIJ71O7LM5bPlMATa0FSRdAqJVDkZVNlA1dG5ihlwvw+ywrDmM8YZJY7akNvw
k3n6VtZtyhztsCEkBGZCsHOufqD/rdtxpKecdAW3klnONO9i+Jyt9uMIPW5rk1E1uxoSKtrDPtHT
J+X0Dtlh6Qa69RAdjD4PV6a66qz0aFxiDWSAZ3RZayvC1rz1GS/JMjmdlMXVzf6KnyF69U9IEBHk
DDLhOm566FhwzLstKfA7+GZ1MLkZ0nx3Cvbq2YB8s1ej9dM4I0xVfXutIlSz9gHWQQ1negO/154y
s0ST7ccvwcmUOLSA7iichF6vNfrOJdySFkEsHD2Y4ysFUpIip+wF1u0Mo3nvBMQ+FfLEUVnFRhs1
D686rowT9yQA7//zhFq7fFRpica2RTL2ROCblIHPJcSlHGwogmFW63kbATRid7mnWsh5n7ZiTbVF
Bsa5dKOMucQaZoSUPqQhw1QODoLznOcdzzQwVjmG3rRCs4dOho4vwhjLt/8bfxPTlEuZyqxlT9W6
GeNrwJ5WijK2J1uvcJA7mp0j6OD2CtepMPY3qn1TrYo5LgtEceBGSMXnbA3HYz2ecmos9M0f5PZn
4KmmYmtEOcy7aVByZOX7J8FMGMo/09vaEAg/Av5lkiyPXFSED8Xez3q4IrtzH6wTlfYR84wOSfjQ
9gr+a+4nq9FQU7jMXz5mInrgz8pFBiaQQ5X41IFptrihvTdDWCN0QtQWioXH0rPNPS4ugPNaQYUt
Pj346u6AEQHpz5PetyqRc7MaVbcvJz2sXIwFvKeMPpdqefgh5Kez3tqm4BaQxdVPVUs1ZYNvW7IF
o3DErN39WFolrevGtewdR+lAM6GHM8aViR3K0gYWhnn2PUBeNeZmtxVchabsxeD1JE7pbdvfpT8F
2HPkPx3gViFD2Jnu6tDjYfpA7FS3Ig0lVjrvz2FCIaZtS+HugBrP7RoaiI5+b2pdhGXvO1H6E7ua
sFF2ygDTDEhaQShkcwUivA4P/sL8HUOgfOdricMKM4l29Kf4fYxyNlKScqnjf8fzjXfJpxRotWrI
5uHNSejNPScw3bVqxLeL7W72Glo4qfX9oAhl9W5Acs1bHiUs5qpFrL34Od0dOTG80clAuu99YRRi
uicKbM56j5bgkic7WUoBeX60ca6evR+g3RDQRUHpHp0/gAD7h8bc+15u4X1OVIve3QxAbFk/V1Gx
vyLVRhEpOQm01pKKPSnURNS/pxNrJ1C7tVFatVqutegMB7mp657mE1nEPQbuhQgU+7KY4F2AX6kv
54lcaHei+OL0NVjBeofngjhntTO4nXhPdt248tIhLiktUwu/8MQdLqIprF0tK2Ou4vKLDNodXWzY
jqudPZ7klUQnGhmJwl1ycU0ZJcFKvw8n2NwGZTFGp813d4KkQquYNsGVTr2A5mt9wcFmwDXX3ana
+8m3A3tRW1gyVyklgLFsnYLh44nBczZxrYPFm2R0bOklwe2IvJCbJ3xM0qppNyNKenK08ntac3ma
ocPTprCjYBPsrlPOMQPbo3IFjOKsawNO5AwsWfr/aYu5y21edcRFIpBOp5z9RFMs110V9KStMSPb
o+L2XC2FkIKZtUH0UsqbmC8Br9NRmQn9V90x1fWU3vPs3XFSmssr0f0k3fe9+TerJdMilMb7F12n
P4RO6Hibld+1AT0jw881gWQMZJYKXQqjgEOw0LX9xtRbd4UJJEOaQQZ9A8yna5F+Omg9LNI0fxGQ
ZeZl3+TwUEyHS0El4Tqoc+7NRwwsWunuRjbzQ4oC/ekcJy38PG3fEiNW4vE+cPUWuKuCq5uVpOtw
4MNmGXoxcLB7irPL1Cq4Vo1XDC5MWuMYSZxFaKPLjfhDYL7FFXjHLEXhrvJvqypV0aCQohOOUYQb
g68hLCmYSwik9hJ6I4/zjrYgOsdYj259tuIpaOgOncBhvwITTaPHsjMIDJdn5MQJesbgb7/M+XK+
uI/Wfh59ALR85Wr8LpUg6szTrcwuTYIFehAhTtn8fBrwip86qE0IroINsNSq5LoKKcZEBnApqjEk
9dN7gQ/07+wk4DNMsuwZolwA5WBOInkPWu3PDrohm4GQJxq216kTRn5XYNCURb1D5FQ1MK/19Eiy
sGyFOYBkzBTyl3/0VVuAld6mTHDW0aB18jOSFc2j+jy2ZtzpkDlP4Nb/CUg1hAfIIM6vJ/+Id4wg
b08xr0vVaGLHaLU6D0GNvVZ+P9GFZl6CYT4sHJzwVKV2hlUbJVLamnj9ycWzLFlmYWQcniD0b1B0
D0nEXNaSP/QUs4RXDnsTABHuW5f7BOqYGW3UrMxBXTwukJSjU47ZFkDI7K7HrIaZsLYaUKlfqERg
w55Kme/MnfaKOzz4us3+cIFlUpYmvGi/0DkZ9zwPuXqk5BexZcpBLwCsjb5wVF98b/1tItC99Ua9
t6StDksySYo8iFwQtWwtSIxRpBd7F+nT8f+xvcvUvQ4wyBHOSAsyNyY9Xy/CMd3dXtSgsuy/Amvw
4D4GhdVGfzRcclsEXdn1S7tgxMEJUzM40Gu8mVSGcRh4rZgPx6QOj4LmU1rDlN+Pdi4LDrP9/Ecv
yf9rmqI8ZN47jmQ3EIAm2XO8/OU18vzjiKjGWQwNfPEGShC5RFxRwxW/pXAjb+7PNErqGkgAPkDC
th5NHPvcTRkeAKjZu4kFz/3eWWnKZtY3P6P0hyzzvvvmzQeofqcTlrAXxjOExyAMUhKGZIs0aGA0
PiWGn5815oh4YKs1K3T3rFctY8jqfgVvAA/LJU3onC7nwtRQrIOqZ9DRCHUX3/+dRaUHhDAtd1uQ
NIlSlIxHA+89nBDEfKDXt96zm80V2RCr7Rq7lYM9p/AY/8GltHkg97p8mWBUUXNhr7AqllMXub8b
yR9Fo1qeqLT18qL/xzwfxCMKgoned2FKi1NsiI4+awbieXDvWHZ1kPhvK7f6BCgAkzrzdgXEgrbD
Qoj2WS5Alrsb3bxX5aNwQM+F89t9yNJEb0HUz4hbgJT2pgVSrrB7fjxJg2M7uuC9tT2xeMjz7H4H
mPf2Eivf40T/KbpfiXVH/AvpL64Smn9H20wy/BA08kC+oqusjasq/Qv0v5GuQ7jhLiOj8AizWu8I
f8UOHmSqYP3ViR8u5EmpzMG7WIrqbU6kpGnHa3+MMGH9vP/GWPRM+Wo8J4SF868sThDtD6wd1S5D
RJoebFtaxDWXHqdKvtMcP1yPTkcVYinRlLdKxXfxG0fB8DEb92XhXW8vxSTcTmaxy3LRI2pWTW9Z
nPr0eg0P//jyJCLzudJKCru4J9i8jpOO4E0RUMkE5qI6WeVN4oP+zOn3It21rCx8IoYpXO+gvsdw
1cmAQ8ovWLw3ekiMOwf94li3somdcluB6+gxrxYp8aLIvCRc7V0nx4cuFuJgWJLWD/DEWtIUygx6
czIRKVKETGudph67wsFGUaXJlfxJ37u3m0LC0Jg52GYxx/kH1GXBVGC+9qUIT2bLgJ9yScFZk0Bh
p5n7sKsXDmI3DbilMIqlWAdEuyrPT5OsUE4pPBBzt28+6hSXBSxaPw+o441ssDT8Jjy8o09DEp67
b9MsEtRd5Am+scj3VCYZ6532HLtmdarsgaEDOs5DT9zYo2ljoJ+uAOaTZx2icfumhtr9QVoTpJlR
VnBqUzanBRvjBM8cojwU2g2mFwBCiJc36mNoe1nK/rQWz8x4xvjXl8qAhCCuRi+Fk9vFwAVtEJOX
VZyH3XSIIJajyJts5/ztlURhnaxV4gIDM/Mv8pGmUQ4b7RN3qVxNei5jqlE+b9NUAStow/9qKnQt
wGDt8lSfaHXUKCD4dbJ7IjMoEYWHm5ouqxuZ75xYcFwxtpEjUgiFEdwmQz3kmcDIgiB7NymHXFBk
EF5HpbOLTpGylNjAkP2T3XaFDoIEbbDtzwhf6tJTXIBAQ2PDJRLGCffvdZGS6yeMoFMOFXJco6MR
obYFxq7rlSH4s3GO26ocon/6RAFaig/Zg5cqmNYgU4JHTmt4tQrwYFIygSFTEImeGY4Ev395GLRT
g5npPa3vt60pofPVj5hUQIamzOQeGgF/KgsRT+6pAVIpzn7Dv6RmVZ6pmn3ZOh8UG7F/7Eu9XDd1
KdHV5UEhW0oVMkWURDYoEbJMgCcJLqRoN0ZqWxqXbmhyGKh2UU/44oETw+uwAXkBxG47hvnMH9v4
61OYahWBZwbMjQKN6Eko/XLRwBkD3zRUp3r+Tp31Xy+1wiU15o7RMnxEs7IwByA1TQ1B7ILm3Lsl
nx5LSfzqlrJvHY0qosn9yUnR7Nr/88H+ahfJGUAyKA7kcSH23BjDclo0rYPU7bEhcX9YoNqMB3A2
NSOvHd4Xqz3T/OiSUYO9FCv7c0ElPgRlusQjlOEoZ9q7xgO9jnKBZ3AtKgu/mUWhjnsUyl5eREKP
mPrKBQC8IcaY+FDCTR5SDEuxE2/lU1LZB1tzzLn6gmYFjaVQeLjkdUlEyMxR4fZkhxkyICrR9WBk
MhO5pPE1kaNu6zBEyxsM7ZGMfX338/qeXs6b4IchtmxHNEtYX798m7/uqEO3xAsE7fs7wAYeDUbC
vJGLGi5vjlnjRwa7P841wTjDbRkzSH6ox3ot1QZy3XEbf02a1son0C3S4njb5XmCRPm1fP9Am45X
OObCER7Eonaizc1MIDezohVfOFiedx9wV0C1YR8sDs3cXwzWFISJ3xgq8CN9LS8uord+JI/Tf8AD
SrGQjJbjKbZJByIubrJBQXcg4i18i51GdcHXPsJevDoyua/tNZePWuX19LmSQnWtraP3wzTZ9Mw1
w86lNvpAtySS8Zk+AsadohGqi98MJKaYpDGrVaKFNhm2tlrTSjMNRXaSbm6RqAgqsUCmaoj9vnED
Fif0S+eDRvO+uPsEoB8xK2VQ34o4wA7rjYf0uUNb7GNSv6L++g/FtCfeu/eBSIcj35u7hVvjs1Ay
tqs5K+E6kwXoKzMuvG92A6nhQ1dF38QgeuVGX6FKS5ukBJ3Z6z6U6Uu1ELIGTz/QAcFX2IKUTEcy
bI/9emvoJVZnH5J8/gufb87frBXCIu89iSABHKbNm/7p7rjm7maQSk6omaC2MGYF9aZSg9Gu2fd/
g2kemPKM0lpiIVHbdGi9PUn+lnecJ6BrvOckFX6gIW3Dy96cvM5Bmn9SpNXliiNld16hWsWL4e39
POay3GVl8rar3ZJGVgaP+GCndc3ZE3l68k4nNbYU889hdV+8S7OWjroGnAw9lifJbCTipJuEBrmY
fx8e8YLMFbIkvKUP2DKM8/vPzrRvkWLk3j42S6Zs+g/TJgyU0fEL9DjHEwBOyrrNV52+JgeiVvhR
sTVfFqCriS+Dii4jkpIF4rkCXU90viT4A4sar8Jk5xftpugLd7d9bPE6LtF0w/A/RBrr0uMyS+Gr
sYlqVmzyqNQSBuU8pWfP1mr8dhRzDT02ngmlVc7z3UImzPbP3mygnNguK2bUqlQoAw84scmxLjz8
T8Z1pYIOP4qWChUXdWpOpIPraGUVq00gpwuNSJHoXsZ5gvy4uiUD9XDRRpb9D1pbMeVXmfRMsM3D
VJxPjw/QsXaC5hcViv7yQgp68bUsCwGxfPYKKm59KUusQ5Z2VTXvOreYMFxlhRCEj2TaVCxvJW7R
yprxscvQu86jcnYgb7lqiz7Urs/IMjL91vp0PWN5nt92LBMtCnN3dp/j3u9MdCEn46ot7sZ8PUWT
jjdBQnChxG/xFlNlRIlTO8+i+ix/S9eGZm//7r6zjGwjmEreR0Kn0avYGibiuV5IMUqibtuSikNE
kOSytgtwa2q9MIgWt8eniPa3u/hbH28v8PHzMpBKRv51J2Uviwl/1F936MHYrN6V4nq4+67XHc5V
MdugHPTnrO3H7AoiU+XGcvT2jWCPTOF263FDZTYdM2DxeaJLZmsLYTtjBFKxH4fmkzLkLYsXjHbS
QCpjgiYKQbmF0uHdMDoeXp9n1dX0Stu4U0KK4ctAnUSbMYIMRk1x5pH+kozYBwODveoG4Tsr2hzc
ls3pVZu1OpeWjoXpu3Lz/Pd1uUaG0WPdQmCltAdIRns5g/044OZqHUHq7BS6NX7W/keTjBYmEodd
Nx6xbX1I9UxSQR2CEQmnzOna4IYPd94a/oWwVBMzWq3KH7+Jr4ZOvgz/cf/3Z6iX87oM+pJdCyQ7
C6i7HEo7gu0aGr4Wv82YHjHgy2rjYiv0+LPK3iKmu0TQyBO9fzjsfDZFlGCeWQ3YYwI6F4x7l0l9
AGUEsu19m0maGMMe4KX7N35H6/A/OTEPca+LV6qBMSDVH4xudzD9MIIdx8C//AyFI6j5YqW1CVLJ
hkJPKz0mPoV70gNIzcHTv4zISlFlHOSrrMxNaD+TL5worKkgPhJyB59fCCNSjvZfE66Q6lZ9fIUn
pL9LrXKduZmdgmKGQYkzCWW0MU/yJ1Wmp4qef25pBbVFt8CR9i9FDv5YEFoQTzE3UX1NTbNfmPMV
iiTbSGrkDwJcad52qw8tZn80Z0SM/oVDTm7GGK+cv7//5opMQq64zf5KNV/CXlNN8EY1CMcsHZX4
wQzApMksDcRk9R7wycHmUiIQnIEa9gr5WuBEGRQqTb+ijqk+PKR00LrTaq3BH8NaHn91L+1a+Xf/
Jr0/RD/skpKzjgDcZYNi76ecrBuCjjLtRbFM6j9x3P7sTxBw22cUM5V9kGP5raCDbuRush8vQZbt
cEeggnQuUad2kq3IjvTBZgeU7DwPPvfzVEYKtyCqW7v3UP5esafuUC0sAI+JRc9DD33MQ1t8gFyK
bcf2X89V6Q2KAsPRiCkzN20i9xgQWZf+6EOT8lNXajpaOXWLhN56vU5Nh2oKS93ntjQ2if/Cg0JG
yr99kq5zPaZdSq7bk9wqlr+tF3uWPlsXXDEwbT2VKjXbEFEN7vkxePorkzVyb58Qt+XMQn+9bBDZ
ThvWU4GrKfIU87l5J+54Z+fEJPwnSVYl9EGfWj0avDrdgImU0Po7fUVR8nLvg8bIZXH/QD7yPlQh
SYvOV7AwZGIeD4ntChTgVeha/zwbYFlTkX9afizrRYqdrRGOu3vtx6XMprm3HIYFfmI9H4QDIQNx
tfk4iXtSFWekLfdDD4XaTULSwHsFOgv8976qmK5fO+q9uEuXx0saC7/uVTL5yz6YUA1sPGdxhz3Y
SHmAwVxyrkXieGOs0omn7K0Sc42nlZYivYMRaXf6Ul+QxTb1YLZMLWf5W3MyplnYHaidrsyBjWDi
k9oov04meZ6QuzYnQoZJO0q90hazNA5uYe+iXzm1Bdj2n43bsu7DsfbtswiBK75BhN+9oNegl8/j
qv/NQ/gBL4HBcNda+4NAxv0rLUIfk3ETfl7CLfJpdxvSBGtOiSArNkg3bsxZa2I1BPIEELLn1ceq
d0CpWjvopuVIMYPEbjvW/46yEmmfdE7C+tJWlAWPgBaUy9F3o+q8AGTjr6bVazVumV11GfwbU3xG
1hE3Gfp44+3xuGORW5iw9GnOIZec2mZ6pOoB7ZyKafvAa7c/Dk7k/vGGN/alAMa1IlCs3u1DuTZc
2O+7m5uNVwKm8a42bw8OupgSC8FwQthhWjcsMcuDOC5NSVh5t3diT2uyjXNI/aVMrPjvWE69nnRb
GdAH+V43GYMj3+2Bjf3FTic4HVqKOhsSQFCVTYtNMHERWHlMMQn72fTQDIzv/K2EpHr7ojXKjGM6
pInsSJNW5WXHZcoxJOblqMHdDF7s77Rj6/6EEGPGWspjhTQ9zf1P2bC0EJTgg2cooGu3ToXccbXg
z7ko66xeRH5y50pwT4RpHXg/DScn3GR8rCJ4VJTXSDiZuR/oQcCkbBXa/IWecaChx4PTnpKPJj7T
GFX6tbis1G0f5+mgiGFI+DGwKoOBYr9rE21k+NNUU+ov/Z+gAdLUSls9yITtUJwvAz9uWtE4G2lU
QQzg68T6LxjkJn2TNcHsEENQaGEOQtfx4va/PnaeyiGZ0sOjpf2dMcOSTyUQPc6/DOtg0J3GpQwn
bvzi/FKM9LQlku5bOn6USV/syTDTpO5OMkVJabgL6gOxOIRngqgE9VrcMs8Hx9ubh09A8imIr0kx
rYTjZnl9Ju4BC0S0z1Wp71ewdVujH6FXcrgv0aSi6sGyLNYFZRkHiHqC5n8RCTVlbkmLTm1OBSO6
c3tJPVqauHTxE/L6eSm7Nsvebc1YMprTPpCyBesM7rlfSH/U42kRN/7Sr0rDTYk/rXr5vt96OxsC
ksvvQyX+uUWFQIXTwVxBIiBO73RRMym2vW5EooBmA/ZiRTePNkbd+P69tt9W4Pk/KGvQboC/Cm/D
1H/b1Oigw1UkyHhhEjYISmVP0fGXJpgY03Y1sjd7PtM/Mf69iLAkVZrtkVerW4Y5xoIOttyi7asG
ZCWKvgp0D+2NzraMv2lVLiKnt/s5pJQ2TRdTTR/3jf793Sp94J+pFymbVvdQwIBk7EXRTdWDLbi5
WLApmwRxY+pB9Ka92nmrmCR8x/r9jCEFC9mDB7vcySR7Zby6CoJV/AA1pg1sF22pQ1/Nxxac0tNb
GAQonI1ZUdMcO9wl+fxg5uZmk1jhVlawtnw/ep/0wUUF+Ve0K/2/aqr36/Ss3NmzZnqVaqOM6yNK
mK8/SloMyQjH3YDlOwJdwKjStukpESo0HW1c37iFbD+fhwn1Yty3tNxBHSuHH+5MfDpVGLaIVq81
F5euwE1l69myhdvifhVQC0s2Gj5PCDIefetd+WdxaLB4Iv/4NIOjeVGSse9rD3DfipieOSZRvKLX
5WL9A26Mr/Dt0mt2mtAElMlCRESIZ/0WDcAVESv30+XwiZf3qiSuUGE5KDcRyp9klczIVsO0lEFL
J9ALKQmiSWUDej9Af+HeN1KU92oDIfaS8FA1I3N7rJDVVoQB3KpwwIxsoAXDJc6lV2Z5yXM1lN4M
Jgcye/bn4mh2Rdtz533gkHpIEXndua878tt5tb7B6iDHDN91rzg9iZITfUrstsHBh+gvYU+f/jOK
Rkh4Xoz6c2srtiftrSPi4b+OU2mYbjAvTvnedQwQ8MCuOq+aD+wwSQHdA6an0/Zcsu9Uj9JZ1F5Y
RVR5f8EQDTrTyFUnzhzgXskoVhoE2e8Rv1pmKBrVmCTbLgu3dhtrkTX2B4qdPZXLF7Wy79UVgQ70
U1E2HM0L92RLphxn02lKln7Jne255QwvavGYOMnoHpJZR/du73u5sYTmMoGX991tZlEBsjEoLtUC
f1TpLKzh+nLJYdwEs0+j1mQMWjdquJwWlLzkOAEqNkHjWMxI+3ETxJfGlhgPEPyO9dRp9o52SK//
gb7iFUaJ58PhYiSzNPtZiaCddEBB21XpLba2+kfA2EY7gWS5af9wH/97KiOlbOd7bRy03mX9t0AN
xf/7bTGbwcMscmPy4L/Hfo9ev+LteXSte+LXZYXzdlqTXCvCLqL/13Kvy1XZoPYxUtdRCQQ/fMpM
mLtiBppCwgPGefDoSDGdzk0+x2EFXRcoYgPtMADeE1hkGxYuTLkNkmLPgq/5XkFe4tM12XNwzOZQ
kPJmKzffVO/LFbr0ZsHy0K1mgKjViPqMCmm3OEPtlX/GbIUk3Kx0C0VJ3gD6YgJSu3dDR+x6qrU6
UkVguzNM/rWPqb4Y9vT3qANFgBwb2tAF5Cc2C9dkwef1Hf6Hy1r2hhUWt1RDED2A+lyvuIQgCQp8
8FJ7KFYQFVRmKemcw91v1E7QIOT41FrnANM1vgw71V9X0X+svLnEkB1QdySaBGIOVPJbudMOca3C
atkLjTr6Xin9/7V0cLVtR1T+h0hoFZfPs7DDNS7TL+TfnlP9XQf0lpHMeIJdyLJyboQtst+Gvnd1
n1CYAxNR1X4QcLTFuLYCEExjagsA3G+1BEUebbXz00B2b0SWcHOlBRaxLk++6WkEHGo56b1lIvdP
dKhqXu1VTRAnTrl0gF7MY1tx4J5bHHJ5VIsNjU2IXIJckGkGPfAErhizy9hl88640gbqIqiuezDT
0JCBFjKW3QEi64wBgOc1+W919LdtMPHftESX+6sQULQ0nX1NyhJhZwiWKRP7bT5Yb63DXPV6xvsL
GhW/0LigEd4VUBpHZ1LuSd6gcn4jHJlqPSWree4vVIG7usCDqsLib6OT3ZOm3m6hD/R0JSBJojeX
F7XvBCJYnwyxSi3welsvd8HxVIIZ8rxU9+NUA7I3UKvORGI/HQh8D1kTzq6keeCfohAfAHECjX7C
WBhlTT+N0zWab7B28TfQprjb+z17nSAnPATGdZCwrNVR/SUY2phSTNcBbt3H9IdTJGWylIvUdEUE
+xObp7BpoELQlZ9+CxFObvt8B1fBlZgEEu4ay8lMKk3vNuJ+GT3mLIylpdBINqtqx8N98k5CfydE
UId2FKTl98w6kMe7sDAJqfzUeWB+xBS+jkpuxPaqjQvfoRQb0V9KCNoiheouiSgka1gC55kSz+hy
fodloMWOiofj/esUlMeP6lGfE9TxoPbF9kzeknL5CoTHJ1lGKkJJea09YnYgo/zjxhnV4yrDZANt
MnoeTRxkH4NrYIiyyeHs4Ilt6Hho7rKrdufsqPxibxQJ1K9dkRVWV6EvjaduXo8drxQ04nSJuwA4
8NoJfc/PBPAL9eUJnK9qpvkLIg4b8poSEcMdXU3EvMQHUvIa878tmJy4dX0LuD8yyYQ+pMw2ZYIh
CJMh+uDMroHI09X6RwtYCBR25JPrpv7PXJTojzXj9PZJKR+UZyyn8ixFT2PM8e+2fzDXuXxk+8xy
gBmKAcpDIdWGR+SA2+pBzp41SBGzErVRRzBPBijxKZzUhZxj4pjBD6i6Z8TBGkFPV7cXDEp1TSYH
wRvBWtmKJNdwMojxx+6y0UQvDu4IO4igaWJHuQS5d/j9MEmEYFfNAk9wQlDoD8ZOXwVxxi12V6wq
GH3cy/nYtHmMi2m6brLVkrIcjzDjKHis2/EcDS5IM9ncy65333yRihhAuYP0s20fDV8ENW2kd183
/WB+ezJZcQXeT2l50veOcS1RgkbHdOzbtivvv6uFvi3+9qs90cCYPTiFLinrBxWtaAYPP0X0eFfj
enXxlhHutDD04wXwQZmP5AtJh3QA6MDkVxTTHgWl7lPQn/j118SaeDcZ47H5rUgKvdpNY0MAXMj8
T1fleHJhL6yQwvb9mo6f83MrO9E+q3Ysu645FtP1iUF1oxbj2Xi/7OqPUEoeka7SJzg87YjEthok
5/r9JePutmITHELX4QTi2L/8TBYhmdYZ9jZoxuUoopatdfiQT9rV/sw/QEZ0l1XDFysrrG0AiNBr
GUUz+zmUXEbR5VGQpfREFUwLTKanQHppjkjBjRhHg1C3sndBu2icCw6t8Tz+vmPDoAlKTw4/r1b1
CHvHiHdxAlIPNm7ibidxd9Cjbjj24LnLwkZohPs/72UUFwRZAefRELvN9yu5zHQodPcI9My6RG8m
pxMLeOaALn4ff0ovg1dF2Wv3BOHlZV+IWXnc6iVzvwcLmCX8mUcOtAPtW4P9ux/fMsIc9M9rLl7U
hAlz19FHw3Fp6A5QvtfvNZsCiSi7ffo1xrIchZcb/L1NhDRiQRWExQCeRTTxsLt2VCOom7sWA6cN
8hZv2Qq3B4jY/yslQjQnNipgtLYz22ddaLHhwljzzr13m5b5py0zjtfZfhLvgKo+lRMkZflyGU2N
MVKnSnC7g655U0yPVsVzmG469hkamV+jMVwIyzq5OXuyY0vYSwHHdWI8p0ou1O5M8GAZUyV1Do8/
+dghmFve3ZmqZk/H7zHQpL8Uq5YI6LD9Vzzvap++M0kp/jvSLQtS0QxupfL84+pSKrD7YkRZHevi
HtZ6zjBGlyKCXVBmk8+4RDGVy2Di2d6nFQsRqMeu9bvf3keY7Big6PuktjryEIfEqtw7bXIfVW39
1+xeV1hx0PNDwZ9xM+mM6UMaGz2pipf1ez5EXdOWzZN1DmHEFNpy6GWbS56mE42EyNc9SQRJBBll
7aYlatU7brSoiNdHE1PgV6bl4Fk1ndPymVpDKa/L+mnCuWDy5Ge/YcUkgN5PIcRT93wp+mckKBRL
zA2AOum5J7d6eD69mKXhC1DYTYcmF+ISFhnX74fUrIeElfbuToTPzi+UxmmG6VcFinV1SHq8A2Ve
MKqdXPeaEvA7cNXbrAO/EIO3WUewlaxy3LVWr+Bk6g89vZhHj/Mp3dFfM3smefjlpLOrNoaO+luI
Wp3z2lmTQSSbKlgv5MisNgSB3URXAo8xO+En2oTEm4JVnj+DWMRq8yk2/58J/SFN53ArqCCUB429
SgEV2hZHuQ/omMnWy8CsvWX3er9w/Zpv20jomnx2lpBaa3wbK5R+vZRyuvIzAwCm35xQTtjtgKPV
hC1ER4EBC1BROZS3I0X+Qgw0XcgMN62wKL1XIveuKbcZVy5CQF+RYkhc/wFtOdfoqPOAScbLV99l
5LDabMnHnuglfkoZeQrQUsAohYSKzmvRPawOpYVqe1gFD1cOzD6NR8z+XfuPsbQrP893l8R1p3UN
1sRXH9ZmJPsUsniltsgX6og06BnNr+Ytwl+d3+892Mtt4k4oexPkIZw95xip+0yo/8mV9XLS3E5T
FGxgR7E7y+OVKqNxCeirOOBKgrSamtURkrTiLkOAIZ0cqTZXyxUZ9TskYJDYb7ggLX3Bf5o2sAWA
Ac6Yu4nv2ch6JKQzXiXk19dcvHeuAILugnFhepBEa8xPf82sOXmjy/Zmp5of3N+25AGJUqA+JeVi
cAlJwY0RmnIyejrV8CuXz625SsjXe3WCX5hJoo1Shp4uRl00GWrRTwEp1XrodZzG4l3YehpIZQwv
Ix63qA2XAZTgUrQTu2FpEvHgld7ivbcZs3AGyPdLz4j1FNZ0N/uJ2r/OdlaYj7AYtaPLUVhMUggm
q5tDh1jKM8VMj404Yir2iZQSz5ecPkZBuGPEpP4Y79TBKkNlKzzDCsjdAqHNunJo+HnXbqACuWKJ
1/OGjO0Szcgutk+y2Q5ZhqPvm2X7Iw+FhYo1o0zF4WqMyqU6g9ZuqmG+IeBz4F5aFocCXlr5W9S6
tty+ENL5OkzXp5mTP8ZX8ofqLKly/ObbRQeX25fRCsbOWykLspe2SkJQSmoZHAHQHX1TDHsaBGBX
+mc2w3RFAGQBQMoUX8fuWDRAEnAmLTC1ykxsezGIgGwKsgoFu4RE6TaCiH+AUWkq6pRT8lw9cEq0
R2Eh5yyGKq2ETWqCu+bjxclDpvjHcO9HV4kbtLYz34ysN+AgJvOYkKa/NF0s4RPj6BniL0ss3Yy+
j6KeI8juoE0KKffOQjAmXSIiNzaRReu5pzPGKAfvKaiiHTBsl/P8FMLlg+7CLozhntdzCXcYo9ld
KzYGej86zRCXtT7HU7yP2xPoJRxDisQGbStKUF8NXZPGjbp29C8iNVtONBSp1uZf30vohBtYNUQB
wzp0uomAV0ia7q1gzNZCKE/Y0TJ4MYPxIH4iz2VFxa8TmPxn30g6PAgu1OxXLpYorkxTZHH/m4bq
LTp5ojezsuZtgtUFyYbjFd62mWoK5ogckWV/5P9SrCYFlXRmo4rRDLDpxKPmuzoKqlf/eGSbCkxX
SFCidDsOrlH43PNkmLYKhc56ByUCcDN4jPD5PEfCSXCyir0gWnAaZGWh7HiqVkYefwRWXDOyG87P
U3U4RPjWEWxHcmS5G8TMw4k4XrcRIRu/IBmDTxY1LAAZYpiA/I29A1Er46dgD3QnoJdxysazBgB5
/vxPoOj073BrcEzH7KqTQr4OCckfkhBBGRsS7gO1hvXIjSRd49SMp1LU7gY/c11nVD2YR/WVHZ/p
YjvwpHGY9iHIG8FbQ1XAOTUhgyKyUgbhBTM0UV5yZoR54zr624rQFPXgeW7B78uyeMKLCXk+qnsZ
K518ULH7OSIv3jm61ats3ab8ahH/qYQ4hIkkFRgDTBWKcQNZNXdM+U1z9SHeLa6TuD7M5lkiaBYp
1/S/GwKWaPueJ16PIzSRR5d9RRKBzFM6t31OT/JaXmhavvC/rCiaXGTxy+RxjbTe4ua69aMSEy9x
LNnt8D6tvb1RIt5jl3pTIVM1CbPz5UyyHyAqJKgo8zYuHDuEXr58cLTzkFrSPUa9y4uFHYbiEE7e
1014uZU2jF2K+Wyfb0XApXAS0E+s+7bZJWUVmuibD7GkHKFQ8BQUpk4dCFYCNt3XxvRTyEa0Cagm
7O9g7RoK/2MQx2eWzDIIY/WGT9PKPil5BQWQZBEqOsVFub7VQdpg5Pq76kgxCRYhht4JB61SVGKd
lEizIVzaXEzadbJINbkLSUCJbaW9MGCygwsY/iM3jBUBAnEsG0c7xdqWSvS2WdGj3VuDCycUU+Z2
ytKkUCaZVBniiufUQDwq22P4QZGZ6R4b5Lqm67KgyGr8ZZGQiRPSwCF+Bkneef0pK/3GgfHA2/7/
UPMRDdkbnc+goA5v76ojXYbvkbgsiZIQZrkJS8vX1C/m0YwgMjzn21n2Er4NFtGAWot5JF+30zrU
/wmTBfJHsByZ3BdJdNExSYdMsKPm7VaPiQ1S/Lxq5+CkD55DiTUQ6vw7cuohcIbYTyxKHWvlu5TH
ZvtBN43H19EN2eNNLS6jNfhrJYTJhcQOdu26ZAZBj6me+zyj9j8YdrPulbwq9nND9ISToBVq8+KI
+U7FmKuXFPxE9smQwndoRKY+iPDjWpVDIvkT0Xws2/6LvxdDAh17RRVylOT2bGYXqcdCbKKzD6iy
xPMAK2Mx7J5mgO474uMovmepoSXE7CnOowR5uIIwORaqCrearu96X3Z+RM9HIq3Gt7bZ1p6toQ1Q
mIQ3zmB+WwdvklqZxdqRzBZCfzabJFjtUHRJwSS/Q2J0JurPy/4aa7ocuYZMTzZydQdoenQqG7BF
ZEVJ0bxfe9Pd4OuJDAQVSLHRPwpU/hCqsXN8D2p+auDqTgYrruO9Quz+NovtDjEFv+qiR1EdiGoO
+8tzq1Ep5FK4Q5kNcMWjOh0QsYdq0usDVEKlH6KBgID6PAkIBHav41ekbARJb82npjR4ZyTPCzeF
kZuTEwCJ6OoRWZecRQhrJqYaXaX5nMOJqe0FLDvRgQ1YMy2pxqdQvDow1u2J7s98siZy0dx6rpRl
O5cogdSODmDKN5ZCPBiLiYH7DLBuAOIH5ZkcD140m4OSH5UDUhmJj9bvD7lVE+x7mdx0K7f3a1Vb
5IwPWSaaz2+WURntkPFI8zupFxh0vojRopo0lXHGlWCzRzZYStPg/yWpC44Y7UEmm+5ect4VRjvM
b6tZoyhYc38uGVrVFXWz2UWL91iMLgSBY6c1T+m26/tNdkFFC69WVZnx+e7ZXc6VEOkxhI0D2pIM
TnKNX9P0estnkq/3my2iiZ6IffmCd8E58D7RDFmWAKTGW+xrd42JBKKrX/gUJUrpaaXyKaidhFOd
+IMq3nMzMkEWilzBMPsNf6GqtFMltEPJNN3DEnQ13rkzTKx6qCMvOsqwLgmQbDGkI8FYETRIrB8F
AOpW2bfNQ8NevXsDP2HyR3bYSRJYdEzv3OgPkkoYEXy2O2tGhPkmOcSl05L3BSXsg6eKbL5xEJJV
JWHBgNlc2rH6PonSiuOf0DBugPOCATNSp3gMi7g7hKg8gRdd1eKRnQrLhf8Su7OL22ftPZiuk/gA
fpi0X6WQ9x1hCSP0lm6jGSe6+n0ZyPWbZp4xlpDD9Wy/SBSbfIZlU6tMBu/7DCge0eseXW+af+JE
bc1E5Axe3bP3ID53UGj+NKGJyaC7wYo3kkmPhFwUPuv2XIo7ZD2YbdaRMu55arUROshJz+KT/C6y
E9apXBe/LsMv1Vdn07O4N/f/FxHSk+BuILgBHQM3cudAvANBwR1nRySAPrriW/jyjpjOhXoU6Fix
A+EB6juAGhbXQe+CGLNuBRKyXNT3o7knFimgQq40UXm4sBEAVYNmaf6xDPLeUpqDVbtLyA4DTnlA
hsDljERWkzXh7dch7/TZhZgv7jEysT96tGuuoufe0gZB9HPzDkI8qRJQpjmXRJlo0sJ07EowGbYB
2L22yzsuyK4R3DkIIprCD06gjiLZ1WHfNGmOonVGvlr3YYbWMTAVlJ4Kz0YvpYJKCoie/1l0Emle
xXjuBjoAl/8re7VlhjW1WSVaM4869DpxoGeBy9UlL5T9AriJwsGMFCapNpqpOqwKG2ZGsI3rb64c
ytNDasV4+8iRWSFPRWQG1BkY9ZiXa5S9u8IWaDRCaDPpQwKZlHdLurreI0/YYK4eya+lZTQU4MxA
jLr0HDPDE3eRZpWnQY/adYZaeMA3t/LxB3aoimTAh1/rFHUiKj1MU1SCNMenWhUlLm+hreb3KI6D
Me4jBVKia3Q4nj5evgbMmpym4BmRzQBH9C+hywtHvuheqhcSPAL/qm5ASJbNu/lBfKlvWckIBJ+o
hEPXU3xwofsJYZGoegvQvHywV7SF1TwCT2rQqYe3w3dFmpRgSvCep3UxqJn6c5h/9jmEkn3+o+pq
ITLqc3tOv/qE0dJU2gmcLHJDwi2D1sMN8g3hxwYa4y/QeIHa6psvJbe01LtLPKcDIeAwIktuTKgD
JO1oB3YiSAozUywmS+EDmkkN7Wm94L2IkqhpsBMvaNJUmfoJ+PsEdZJSfdCsrlInjcm7P0+iq3l2
M0KKyWSa3s1L9u3ZjIzOtBK9s9SCOJBs9Wl/FkoAJLInNZCkE1Dmo943MMqNdAPAYlBvXQDtd4In
kj/CR4ERW0wcKkJ73/1N3irxt2zIUGy4WcsLAloK82X+OCadgtnR13cFz/9MGka3Q3quqL5cdhKi
decsZNkeIXNV4oZ0+h/YSSBGaOqbE9jHtBk5nEE51JzvcuB1mTqvPRxrHfBBl8mCu0Xdds8zTwlT
kv6mKY58lYZltXt2ItcNWFZST2HYtVM7F/TDC3AYdlcNIj7wkDWJbu1WHLT7WQS3A0khrx4ytbIO
q97spn3+GVCmzvB6CUm0SxXQXz5sEinEuN3x27jkVfQAm8SpOFLm/vWm7xYRBoTqwv9WHy8AbESX
Z5NfE0m8WT+3CHOHGZhzF5hCSOEcY/Nj0lt8xSq5hnHdmLKjCD9YFpaHv0ixtCJmiUB0Zuhxnmfh
AarSrExxbrGzZ35FJcrMob+Qemsq+qSHQDpEpaNqAXaeFWHP+HJRmFbGoj2Z3dwUxRplFEnOhDL6
9uTs75X6Agjk9c1xrKamL/9fw4jWZfEgSBXdqr3Cy9nRj+rJxLBOhZp2jCsQuOUWIznRtWfjcdyN
PVREKveEwlAg8bZc0q5ZTpDs3CgyQcjsnx+Gac9c7UmU9dwScIIKsdro7G3RP5sovDvnKT7QLQ4W
CYL726/j1YTZ/HufiAjJQhOqSadGHAj0BtWhfbKLuMPcfUwpRmT14bz5l1qAD7GWw1hXH/myUOSN
4ALfVQk1UvLRivvfB89yIj2hFBDCld7913UR3gBiG6V/MhLj8EYNZp1wITmCnWNGXvQQIK1V2D6c
q2+Ik0ojeENNnACPPICo5qHO96Vs2n1PNUoVaRAH/4bFGQFCHC84kdTHjJdLxww47SPkr2l6tVqJ
m2Isr/I/oP9dlUc/lpH8OCSZhEBhY9X9GwiTXdLBGqWaNeZk2EbR+9WhU5j81hdYdUkDoVPrFDYB
MUbxjGZKFcq8MqqiYR/xjqbEM3tvF2WwW0CDyT+ghTFaxtw/KLDm7618mCd+KOQB4GO4zkp4WQ4T
+HVWbGscyU9fB95mKaeUMk+vcqtRKTyz101dZD7G/B+Jq2hK+GqRl5pqYAqs/wnC05t+zK71Tsdd
IwcuJTEKSmFBOShwHL6k+Lp+nLn+Zsxrjpv4WuQerPss9P8/9vpz36rxBO9/SdYYHhX0aKbQVfcY
4GNultZFMxfkcV9mu3I0Uewcq1R9/FiCzrrVOH7JfDtQ09lT6ZiL48rufX/I94rns2OJkTu+0fKl
vu4rYzKSJQQ6QaHpaVomFpfeMYq9h3L0XCjcvgx70pmCroHLPCKoYIO7TgCNxMey5rL1aas2aFU4
tltEX4nw0QdTnn1p1SdUvAPusYGm6ReGXRTI+B0pwVMEt8FgX9V70/8MYmx7YegR2oPsSl4QiJWS
1klFNrg8m9UOSv+CboUcMwNmxghiYgF7WDk0UtjDp3Ssf/5o4BVAyX0p8SsSDLR7KYb4FSmsxJ46
bJsaOXcC1uWbs/qh+9UU3IUhIrCs0JGpzyj4+x+wKHFkqtR2gCpJzP01CyPOXvEhWqQdD2qwwGXZ
8PAdprxRC0wOgPy0mA79fIUzMVdL+zlnfXaFQOOjfYYeDGYtDz7Pq/gQgqDoHqyYDQfaTUhb6qJX
faqeRml4ZaBHuJ+KSJzuMKE3iWdsywqUZ11huAbWFAoTmkqEW/s02Pv3yXJGRNzCsmvknhdleO6B
nGwOM9Q8qgmptZ165WDopgwNuL5zAWlpcBfBttfgzPiAHOgWgDt0uDC7Isua+YLV+S+PNE71tCWm
HZ85shYtqVz098ZDGZrBu/4ZgQqV8ezm8R0+Zr/10a0xghR0WKh0Vo4WOmTKBeNFzXEkA8828btY
N4I60MA6ifIKLEtWkV3ALkHaBAu2F/4d9+/3oDIkhXdtqITnWSsp04SIQlzn5D2Sh0oVPEI+Z0g2
kboYmuCCGsDbv81pzOwfjgJmmRiVTM5ErRvn5dEpaisAGyW3u7eAqBvu1IRHlHv2rpOjAfnjgoBz
EhUkQ3N+rf53K4IQB7/5pdRMWROaeX7x5DiAvdV8lhAoUxf+ZCjZs0/dbTlyb4QqVVM2tVICFr21
ObcSTzdtIc32jISV7pijcSSyeg71EuN4yHcMkTsLgZjrSF+wqs7h4D5Tf1/frk9iJEMDOXHloncO
efhyhlvtuoI37cXT+chBidPrvlUuMklsPnGZuk99LTfNUigPMl7CWTB9J43eW9GWL/mzBqtmuoDh
ORHLI7xEYBWw6eDLByxPN3Pqy3+B264v0/y6cfsEkvkMlHUazOwj4qx/Dswwq1RT77Q01IsSTZXQ
9DzWsS+9pksgqWGT7g9MwntOG8CK0DlH6ujpHG234XuazwTohNPmZM0vd8fNrbETX9ulajQj693G
mPfzPmTY4nojoOHBIjmJJSeBxeG5M3HPYA8yZkngFTi95lOKmrtAXSJXk+Th7+HvqeScT/6aWaXf
DNIAPIzx7cfCoWNrtrC9p+oc1rd7TXtK0KOKA3Zwq91Ky5CAxzx8SFwLMbV+F08gEHVHA2PghIdR
FKdtZ77LYaBHuHo3UX0/gw9fZfNdOi9cW+dozDmrpUH5jSkXqRCTVqs9D9rKM0zeGcUVM9p8FKbO
yZxZ8sujBbROAhUajKIWwhhxKCV9Ga7j6Kd2tPyJd8Y9OcLfzjoMi+7RkugpyGykBg9+mPwP1bGz
YYOG9VXxbf9jTAXnBosyqj0rcwWNOYurbXe4oGfoqf9azwIyffk+v0qoRsTy0WmR90UcUi6tuTV9
7Ng3C/eTzjtOo6YjNgFU/t9cebDZp/lLM8RA+Qy3AbTNVvlv1YAMc0sA3IH6u3KtzDoUhpx2MFt/
kp1vGnZCbDUWDRnIuHNsAJiEnUaJ2dyjQ8N6E937fwAZoHs1zKjsESpwMTOtdx2+ytkIRg1L2W5O
iy4CTyJByUS8sBh3TjV315UQg7b312zFL2fCHmfzoxJjKnp09Aatft5wbNYaT2an6pBNkyB250Hr
sHhVFTAh2nU1Tfivvb66QWUHQiSrLW1FA4iVAFrKp9GFwsZQiWKPnQTMrw1XebUR44pitqFq1H24
VxASyZIFlUsY4X+kzUZcxxxxRwZmgf6j50Xp8qo3YzKc0nbzrICzf0s06nJQ2adJJbalP48CZt7Q
IzeHPgwELp+KbAizfLQ+vspMD+EhfcrPmGbRkNk4cH4G1rq9JV7Ip38KBhHgV1pa2gf444aw5uzA
KUsO0vgtc2mCro+Ui20zeN4x5OdluISqtFKiXY6J30YlfpCLPOz5nimRExCj9D3ldSck0u14+wsB
0Fw61zttZrg0DCPPJzcjAkyHQmm58kNTQoCZndguMm2wKEFoZFn/hu13+whZ+5qDYT5kG7DahCQb
9uNwCTGZS8Vtv9lVx5cibLgh80SdZRaY1XnbVwquj/3l/LAprGGkNcQ5J8LiY1etlQDPelsHNPP+
d7PtuTQYD6aJ78A3+rBwnDfu4b3032U6vv1UH046wIBpQnNLOG3V4AcRJRojg7SwtUQWyiM9A1KR
8gZnwbxidewPmJuc1RCx+dFlfJ0/AO6hU+C8qexfi0ByejCxSqbG/GBP56mZS1dGlf2nucACfxq0
W/0tZPLzRJ8GU15Y8MG4wvrRU0hlM8SAdfETdo0vdE0cV1Nu8sdo4Tr7wryPGSsxFUWQLp4ehxfD
k26AhC65qohhiOcm/b7uvSVoAv5I87nkQM+1wQfF5jzsgxGjCgJ0R4Xm28bTMUSZlqklvwvEBsCy
U1+ztxlb8Tnmp/GDv76uj/DW904ApIenka+FMOyODZ10Ypj0MM75Z7nZrrD043f7U5fvptpf7Pum
WUpNa0kuXrsgPO0wSv7bVilXLeTrb2xiN6tSmm9loD5BTyrkTUsgLx+JxDDa1OW7jtNfcQpgcVuR
6ZNmjnaUXNfyubhz1hUixFDP00Trk0yCJk4durCqUG+KP5dfexVgx2VsjGGEsF18UKpJLsZ+j8O2
q4cH9yqNoVlT+pCt+O02uP0M72KFdlIPpECbHte73zJbNRT0DTFgnwx5SmEexBWeMaceNlKO93hM
GCrkHG/iR0uFwztyMMqzCunpky/QlvVYDlAWZckIDyYiX7yEqa7B+YDgvOsTSdSanRy13KJwgy1d
IdeJUrfYtpcr1hNuUaaxm46mdjgxcB1z6bOuNZ/ubFS5LeMoUgsM/HzPjEQd5AMytITNjbb/3ysf
vT+0+nYs0rMVfi5vCs67hwC3L1r8/mrayDmwcU6MWQcNZ+RII4k1wPV14hbpJzWEGPQSoV6a+sQ6
ND8G1GV/aSBIEqzPYcZCo2BOb3cZ7KLrfT7hJNDBClh81Olukn770vj3IKzAMduhM/wFPxvxhSts
26yQc687V1ga9wCwWS8h42Y/vQ4pvf8kiJvZQVBxpxmX9u4y5xF3vnf7x523605DvstF/7SmjyJ2
aXg9lMEtSv5XOnQvR7VV4p1Igjsbk6RH17CweCf+TjsWtdztY2wT1yRSRZs31wWLXbZQlLMF2lA1
Rc1cPTFAyBwAJZBoTBCOUhZ8xrhT0jEi/XlX8+TcxBgE+gAUSr8YCY8rwwVUxFn1YkgL2dXRF59O
jHzn+3YKKzahefpmYXMH1NeR4ADp9cRA1AlvZq0anyoB7KbDHj4G/X8myFsx/5BHiqbJv5VBlJgL
qyB0tBYYF5uB6CY+EWt/cvSg1rRO1BcDmaaIkVjImP1s4fqrznt5k6hCnUNYKE5qiN+x/3dPcq4i
1Sy00wGl3t+TgOThd1esTOr1n+5yn+sYxS52GITpFsyUoGMG4KQ5Itg5TWE7MrCGaBFt503p1v6Q
k6xcbLJHOv+vr7FOCJEHxLLaodaM5HmTxrScA0n/k00D1yTxGyTB4Nw9gST62qqktua2ju4/3KFp
ET+PNuMKr1MEFw3BnvW2Y5sdSO9zqz/5ZAiSDkV96d9JIveJr0Lq7rk14nTqsqW/v8bAq3gyB8ku
FjA6+vNIjlixtWT/VHECAOa8TDE3det04uA2bhMa3Zj0zcHMOzfWGHdhmh8bLhrU/sShQUOfJBjA
vNdzxUuOi4eL0BhTIipKzMF6iD515G4dXmpu6e7veb8h7mUSJ6xutxKVHYcaez9FoGx9jUzagORU
iclfnpNSTGI9lDoV8fM7o5KulUz+GnmNX3yODe4XvkLN+1kyq3a7aOE7ePJg43IaL4ioTjHqaSFC
T0uehrF/6Yym4/bTDUSAYDpG1j4l5/y9uavQmtyNNAxDizJ8yFuebwfPF0Dp2I3sagC5IsEH9VBZ
78iQNJFI6xilYmr4a9ELB0xVBWb6xbNQhRTMcLD9KxgJmtdD7UiO0RUwtWn5XHqwsNEmIm6BkdTw
JJWH8wyWDlqRlL4jCrfRhTjvb5RdmqqWcZStz2TKmOH8yX8JKdzrsw/hS4kR1slVEZu35OheKx86
v7FQKwpwUsvLfWtOiLQuBnSvjJGnSHp6Aevw/RYwfWK3tRbU1zKmPdJrtk1UtQTT4o3qgq/m5M6e
nVuu2ePomuziTlRncv9JKQ8ETSDVm1uIYrCMWmayoqqSbYgA2h5XSsPCvEJ2Mfo3dRcslGE3x/dr
DfhoL42OlyuHkGPDQXF2Tf7CjhD+SBQozdjlvviIrT0Wlbh6cUoN2JdIM94abXgTNdh0hHk55lar
1B6n4+Z8EkgnESLOlCNWG4TCkXOINw8YJRyotjdoWdhhuBavD9YK7iTfMzK8GD7TfY0dhgDE6IqF
ttnP9shwcoFD0jWTh6U1v6T4+TmzNuHiXInGRIWKEIxipbOw0UAknq9xFCfrzIj0GNNMiNMs0pJj
fYs4e9P2ZZ2nN18ykxIhG8ar3nfC9cb4XQ1RPvo7Ybu1KrDossfCTmgCDrabaqPPlMFEvqoLwKHF
D2ipy+Japb6umFaK0pyCIfRDmODO7G2tXvJvTRuwVD27Oj/MfMYclU+DgH5H73t9qDri6fEeqpss
4a7nHq5D5NZhMRRD/LjKR7WpOJUVl6wfxW4bKJigBXxIQtbxJe9/Vv4n4zCvuRuoIybVKrVE97PZ
THUOk3lOe91bfXvzXiwu87PuXupyU4qHQsRbvNtyCy/5a0rLUshxkWIpmqFHydQerhvtuhT6MOZS
Ce7lj2sjEfw05igG7O4ePbjmInU6CpVGf2ON87Ye/2Tj2Xj4haFx0t5eGnkKxiC4cWTOMyzhq2Ez
LwPPOePWMEy8rH3YJRB/ay43VnmtrpPtaSXep8MTjFx29vuqjIO6giOyjMf6CmzS78AT/BOX3Veo
2eMhNBz05wGUEO7eMIfqVdpyP0HNA41Y2GO70Htu1NX2BXZ0w2CROzjGfIpvu97rYHxtzol5x4Lq
MR/lN9/fdLSggldf2WEZBtrM/1m73HCEmn9MSmS4RDTE0cSNECBude9kNU+qAsmAZSj9mT+bVKDo
n6iKEe4wdcOCdZnJFkHnNdtHMmQ57jIV47oGMqDx8CK3di3f9rMQOGchEKdTzffscHz6gmqQtp2K
Dk3KCGF3CltKqniOgqjDvwpFVWtbjy4/sQubmDbC3bfqsJxQKUJz+bQLr3vFF3dumnMek7XbKxIx
/kn/6yecalWH131kg0Wcug7N35BWxU9HkQE4qYZChiz/ESyzbDtwTMEyZKQtYnsceRllvSLoLlha
khXJMB6oWlne7I/ar7vDlJXTMWGFGU1WqJKK8MxaxsAtHWHz+m7vAVHSznSntWTuR/7GVXP87YaP
qrnG7WOtUehR/EFCRWI7coH7fAJXVGXEmw9EEeP7xswa7XqwhzNvKzsv2XLum1m9dyeE2K/J3BRG
heLRAo8+STx+LTI0lwmv1K7YN+Yl8v1cEUi0qJdzr3qze2sBdK7GaOc4sUaZ8hn661wfFTo9FWHD
qxEPEiVQ9PQ/IHTn2QZViD3blBiTUtQkYf4BPQe+8Eo6Q4ksiNdqr8yB91PsVXqx1tUwu61EXZCH
3y6he/KinJ6LcP/7qa92V8zNoJ63/x3DeN+HHMuU/cfC76GVMSvkKkHMProvtAJ1S3zum0InUW1w
5dJp2DYNvOYXI+DCrxqUiSyUoWeQIRh74cjdBnENhBhr9ZKegHdHxGNUp7/zCBuUvZUJv3TRxMcJ
Z0MvG3edTgw4jn6mwnCEMpi7K7XWX+PX6Ap4v0PC62yyeQa/17vLfW76ww8KevOrpxE0FdAwOd20
XQpF0zjtpqhVxUwdjMMYUznWlVyIj+PFNIlOl8Q72fM7uo6PTkCQqJqROf8soiY7mGXf4V1vTAYf
nso60f93pG//xb+V1CyY6LvC0+9QcBv9qNUXxUs1KsdaZsHmWie8SRa/tR98ScO7LI43Ef8KSYgA
Uj7ITGL8zhdl41Hl0SIwKG18Dab/U33hXVwhd7AyOT3/6e1xCoLk9b3lVhJ9N92GHUXKQFSxD5tr
kfvIJ08/FO2y7VqgB/Kke/G/XxlxBrLsyPJeN0ShOZMXPWpo6Ty5BsVRJ/8fM6lASxiuYD1ZyfAB
ufzjecLHsiNI16IW3LDeOlCEaH01u5U3UWSZLjdUGRmLkX+xWYKNQopuEusYH4sO+3FOH74sZGvh
B1huSBczI1WZvo87DmMGVPJ3fc4UEa/NJzs3zHa4IhGIV2CI4Zifz2H4EOm+Dj6PaYVLnNtoFKUv
UM0loWzYVCj69HOrkjXH8/HhJrIjKyYADEO3Isoc178ridBlQqr/sEBK0Wd+A2/IiA/W0ayNACXS
lplTfFzT3YHXahMTAPVqYe9vhwNNfaZZESpbsAW8oPNedrKFTuUG2Aun0PFOMWz25CTe4Y2kjMuB
cwNbtjUDJVtz3z2Vvg4/5t2zdE5PDjsji7YzHnR9UjF6ozaKzWX2DGjSKLJF/MW2YMFR9vxYJv+Y
o/vu2/aVNGkZZZZ8ZF2esQ55YP1ifPaOrudeIIhKHiMaggI/ceilCfVMJg7RZcyDdFrzgUePeEPm
ynJ7Hkjr0GC2tfWJ5dFJ02h+Fgb/GXmwxWhdavq0DAzfIjEN7QXak+u77IIkN1g5biVovYyEo5Og
Lp65OV0cObZIl8ApIL9Unhl7tAM5G5zoFczaVZU62lq8tRLGut3HwFy3qWMscAAnq2uUQCN4hc1Y
KUUe1ViZ9i4ZBxUrtZZGctk8qlvk8ky/RKxQfDOZydlw5JGXxGCjnvxBfV7mWJPAgTpbUswl3+f5
zmlJ7SDkerRSIbwE1EIZyjuLI3QYTAmjQIdI7j/d6wgi9+mkfGYa6aIJcOezeIxj1m8PBCNugyw2
Kuo7vu97T1tApq7MVlnKVYovoTj4WDCq3gfydmWhmv1olemxEvgV6t7Rw37RzI6rC/c/V7dUJv5r
xkSRxIjUQ5ZLrDwVjZ1zWsN4XfxT7TZFP21Tu7ymyIeDCmh/6jLjE7Fz9Wa5uNDmKcPs0RWI7hDo
rtHUW68JE4CKg+5MC2yDgerIX5erzuBD1ApSBJ8kSe9Ge9YHTkfoO6RdHu9EArAXdprFNtw8hDDD
Ldd8J5ScIADq32+6zIId1zGlMKNrp8C1/w/E22GeI9ClvtBghVlEdezkofridYhQFF6Flc3XBEn5
TX7jd+jk/7y8gzLiOZ3n6pQizS4T2x+6E/BW7/6ZGyhCjQp7vIrpfikT+ZyowG+goAOFXzQHGUDv
0U11uDozWW5bHrfBH258bTWJ9ieRvbONkN4F0sM1QesGNFb/V3kXcATpUyVoJGr81sl91CpTG4k5
l1/uR+oHTtMPQUsZzAot/cn3MylA4pGUD8LOjNDPBUYlC4YfyXVctOULCiMb/2ZJiNrRjGBXdosY
YF1cA/ona21aleQ5DPrkLGBABpAcAjrD6MjlDjN9szvuOC6zGJHW39sGOjodBQdYFWmxNz7pJ4n2
5g73dq/LUr6f/zdRbjyKqSJ+JORx1S5x7wnlt+7/aKMKUborTXCDT/mQ73wLXS9j6hJw/YucedFl
M/wPwn7RaxZKfCFjDAt2Wx4Zprq+8OWJqvrqEztv0xzcrZrSMFpmXjjkrc2fVWEH9Vh9oGPcbicc
KfcZ1tHaKtNsv/ZRaTjPuoiSZOReURBwSLpAUOyoASJeLtuGjQCnEmMGfFQXYsqfGvpb5GmODi2u
Dd4xZvkrEzw9Fhkl08fXBaNjG/1nLOwObOMyfXzrwGdHamjxFK21xBo7lD1nolrGHY9D4txx5Enx
kQCP2EvPrsbPXTYPHEpX/q/lDlrITukuFI1haIfBbAXbG40VGrLdydf1Txah710y7X7ktn0mpIpi
/FQ3zMJM8w71lMvntexN/xJ/BGrVj51aDaVxdhzF73QfRXp6S8Ejr5ToEHvnyk/CqS9pVyon92fM
m/tZO+wir3BKH4J7OHmwyfXwOnS2dktx40PHVu8w936FsTKLCGp7wjKXqE+p4cEUNJ9fgH3lKvle
fWoTCQFzabn+7G3vAaaAMgRw+MGlx/7C32t7vf7EvMTwDe/fwQytnFyiBdTeu0w/La+cdCbENbg1
UtHcLAZ2uY9mro0hzHDxh9eOxlNLVPjeScGvxWzgXo1c+kgLYR6XRxwj+vBjp5i3JU6hl27aFxrx
YKLu4nkdcND/PLsdun20bt5/7H1umPUiI8qtDyCzWOwhOQJAft9ajvl3dK89pnsQ658eS/jpsPtl
8oPjlSjuBaRPazTnMik8PF1CU5C7oNtJ0IeMkDCcJx6fj1U0vSSRQd0JEkTKPjOXoLDLIR796FN/
sezbOJoI/DFeALLmCBwnmnxPbzDKdWOsTk1S7tx35VAmu2RjqZA+KwqO4NUZIOqRcaXr5K80hzSH
dmQjNqz66BUKpthIQlUPN0XB9lc/8W5NYgjfXVGpH/mDCiP9RcEY8UOqQ6io0dx/pmfPVHzh5ptn
OjeNb4LtoPDc6loLbZAmuW26s3mt7GmSmMb1HYlfe9z/vBWDMQd99i7HEIx+ap3YQsjXH7oVmvea
lGBi3byxNzBNF13de34xEE6ws4xaMSFdAaiV0l9rK/WZwjSNbrw+aSG2+VD+s0fzn1NUSUl/mHsm
ukLDRZ1uBkSo1fqrk3ZVx1ixwDYjssO1WftoksrlFa8WxEWTa/0h2CVGcYAqtmsiAzfBRwl9vYgt
98xWUTm4KaokWhhGJKrW3CbvB8blmEKGo8xMrQTLfIC+tNNa1JUQ3NyccWlPxRaawfrpJbhRDPPu
yKtwFgGBjmQaUsU4ooUVOFCQZQTIF2VTR/9cEom135ZD2/Wfj0j02/iOaP4dJe1lG1jIN9yhQY5i
CY7jIKU3wFSymDwDlfyfNS8QxovPQJQGt2wqZh+g2ZLdUY/Am3ybALWu10G4TZWGU7Auh2P7R2jT
3Nz/jNq8L9hQRk12OqXR6N7AZEGOa82JehAcWSd085r+f5HKOaNtAMTsG35qRtymIvU6Jb5blvw6
3GfDLL+8yeW/7I33ucesMPcERnQyt+r9SOCk96QrMqt6JpKDHWBhZ7KMAu6cY/tlLd6uSpbz25qx
E49lPQzoqMTyKCbUnY92KywPWtQe6QlkgqMMU76XhT9RfiNxt7UHKmR/zTrCchwQNDO/utFzpNrl
EDo/I0WsTMHOsbiIzefkGyi4thOwy+6uTr75uQ635ygOE68ANhs38tr6k123wpqXk+tnaJb5XvIi
E1kWmXquhVVlil+QtX7CHmJYhOl5l8C7xxx2qfrt93lqVZv37LtblONQiNUcfVx+i0sJg8vO4xpu
hbUFVPX1TxwSc2anE7s3lrIHNl0O8lM+r+uT2MK0Pe6SxgJfO03H6F3qCiQT4iW4o9ZCHu3/+eP5
E/DXABHmAhI7sRZSbkXeaqibWwAXY1iMk6O1MVig9K0RdS1EMOxlxgIqyRQKsadwGJ8/jr5unDJP
Igisy7IlqtHbtJKBxDaEsFOu59hulqpWJRxKYmEOxqu0hGeJMe36uYVZBOPC5ySQgD51iGxd7glH
RXNa8Y5mcDsXapCGwo2sj+H6FnDZBshD4QQPbqjY6yd1oBCIl1YhvSz2FJzUuc0+izjguytou2FH
qXtAnRXKa03/RZJ9do+36LRvuMaQY0w00P6FFBk7ptSKYkkuXk5G3vHwTzugna/29GhrQ3VgjMVl
pqEO3BYGevojzoOaqLK4e+TOB+MWVbIVkRv1++SxJaAa61/ceXh7XhF/AwrsglnMFuobQ/Zj16mn
V0ggkpb+k0Btz8egRpH9tcc/I9wjHbca1sWoXxFawUrRCkPCDlpbQOQoydn8It7rdsPjo4GtevaQ
jY8IZmk8qQFSftZAPEXBcbIRJGpJ24sGDmliCtTAFATqyL9eZ7q0zgLebzT2g5lsEorHVMxYFxZp
s33qBELc7f3SbC+xWfi+ehYYIi1yHMMso/Qd9yV+6lDxyudiDW2qzwPLx/anVtmqtiVx6eqD32O1
r4f79NJ7bCFKsRJr6DHsMJpw4T9NcM55g32nHbmYoD6spyExxGkMZP5YOkF6VCMsibRzsFHdo0co
fMvm/ulD0xww/jQdNIXOPccyn2FaQRAJ754ADOAt0Rnn+DXRRhI5GAkQVP1h61afpi5PfYd4a8V1
lxPXpPSeKZFvRNCfAiWR/xdmYJ9kfR3ov4Qf9qlSTZPDWeZSYFElyUFmy68QkPxySLHl7m/tQ7I3
WQUvvMBcuOvxBcjZ9VOjcuy2XRS48LTjQWMWkBIcdyfuIFrtFU10cAoNeHzoq2NhGO1YJozRn28D
+fZAzFpFTwST8dbPBXzDG1GHmV3o2JQXZMALY04c7s0gHCOOxPVVjQgXMq/A+xe3p/OJq/liKM51
xpf9yo/G+xgZGNGWu6RTaQxuww2UgFWVrGpQg8GdZtDJqyP5lXblmFwnHK4nTfovSBnQQGCcCd6R
jvdIReOt6dND024TFvEPmiKDMuIYpcem+Wn9pSuCPd4SJFpLQxZANtemaLoJfqllS/l4UDuTdNmb
R6DmpF7E5xAT7npzIsCHNZ9zRFaov7Wug1nG/gdVmJDi2DlZVv97mLjHjYh+hO4JRnlSUXX4Abpu
myreEd4YXhnHNwfon3ZuYYRVWEOXEjgsLB+f+RAXZoK+40bbnHjG8nOQeQxpH9sEOXTuKbm6wFmA
sploK5HEruwrUF2s+b9h3HEl+Vj50YuVweNeuKoycWnd2y2c7GlO2XUDMhhgUvmXeAjec5aW/V5P
TSlUG6opFQjimBjEDX7DfiTVve0DENl7yVo+vq0tlRLKuXuVqZajls9rxj21xSZMPPlqTXEuBnL0
FvImbeZR1Zykd1n2u5U3P2PJn9eXPBI68swIY8ib3ByC7MzFvqloLZft+JOVad1NcD6OZl1Pt2+S
ehZqjojGC9JlyW/WcGo9BG+vXepjJdCS7mqixRibZle2usJyahdm9BrX1HmnutUTNM43fbK5cJId
7Qh5MXUmBK2wkg7oh2x85kVY1BiKUFJUajgBwzdcXxFn+cocXPgHsxFLVVA3szuDCZxvAnM2an6y
nRp5Ay4of3P70G18YJaMjVqnvfEOYOHBuokWxk9NCgQChidwxgryXFp2vCbyg4v9f75mnzN11bsA
pWAowXMqxbxbNWTmiv26/XlGKlvEUPqxcJU5j0M5FA9EE5hWc0Jl3tIht2Pco4mcS7Z+J+/1mQWa
Gl94mJaROx7UGf+uOpqnjQCVUHQ1NOq54sMxcTA+6o9ktfSnpNVYQSkekJGrs/VnKTxGSdY+HvbR
W7m2aNe9V1Trym8M9KwP5G7cfMZmXkFyyTHB4mlxfNp4kCQ9qflfXdju9EMUCq5O2MkgydMccHeo
G/JuwVUp36NH4j/mSw+td/zIhgOgiLcUVmzNHXmcf5I8ONHNBqgldz4iVH0miwWPPb5BhzdUB734
VHQq40Pd9TugVp4HySYWAa1BRRyXJbIIeLKB1B0XU1tAztlfGKmeBVPBnlxnkOsS89JsImJMPpWR
DrpgrSpa4cq5WQo8fFJ3AKxaxp5W6a1U6aJeFTcStd1OraRw3YriKEVgMLi1FrwlqLK44GwHRSG0
JDXSjy5ZNIjbk8UJK3EJu+zOIGG3DTy+K1REesuNOb709XHyUYi6myFMKsNPXLGTT5XAWpV5Gf0z
AvzBJEOJmTaGIW/zcxn2rr5G5Io3s9RoCBDIdPJMtKHA5uqEcJBVlOTFfy18ZAQrLRzDEgJwDSDQ
g8T7p+KqCuG7xn24nQkLW3vZREIlvXMPi5rlu+aR5BQHpdA+dVswSD1yeDjG6abaMBUv3nNKAL+A
y75htOLoRyEP5qtLcR6p5KGc9Jr9zD91JYvkPr238R8jOjUGklFhUbPMV6xJNdGONw0gj74EgDW2
y3tNHf85hiF9DVxWXwFvMJn+waDyifkZk24C21C1rxw30wXSX+MtPREOeSL2lQ0KAdvmC9R/3vsL
/gx6nTbrH1WRtOZ0s1onuGnlmWO70nXBiveMsmiu7qKKNmRHR4pgOizLjriF2F0f6pjWJaaQIn0X
CoaAYbKbL0KiqvLQYljaR7tMN5OszWCpZys3rlED1PZBjnY1TsPNJ35Ha8UQcg6SrK6RVmdBgUqU
PN+D8R73/s/oyjkE2MAm++lEKmvnqH4RRJPrtN9t9ln/3EntbJl24t/PMKpEK4erS0VfATVzYzFd
txw0rG5lQ0JyVn2Hy+Hb/k2c0knveFM3CXs+FIrl8ikR+mn7eS2X0WjxovZcODBLUQohivC6LDrg
O90aLGdqp8JVL3nENjyG75zUIrnrJ6vYGLU6HWMA/YSA5V/UXouQG3lz67aBCvEMvYRYC4KQQMc6
QJ/ICcE2siiWxO1MCVylUNvlBT2vwCoFcaAh68LM7cnd3l8+9aqAO0Vu+Iq8W1wgVMZehVyhWHyO
HalKUXyUEv6PKhAF4SrbIrk96Aq54cnK3yGuV+lDb/r/uw0Pw6Oq8RdqReCRtSlwFrTnIc2ojfxy
WsvZxIuYvyd5LCITv+5l8eRMxh/axdaO6sM3oTH0K6Un0p6P/vwGq3HMvRAhLCOVjWch6ykDQtG8
XQYNGbx0B2HJ5kaxw/FsslvUrH1Xe0+800H4GYJkEpJ/8L/4h1XZUx65XicM+Bh0bROp6aifaUpt
qq6gXcU5PgLThmyDJUA7xraUMlHwtIujjdjTHJQgrHOn9G6KJkvQ9XCgN4VVMQrwqbG9tDEggpxN
K+6+zQ9Qsws8NhhLkAJNvs3EY4+eVsk8KWPQDNRN9ufoD38f5+QKxf6AqZuq1xubnfzl/42DfiAJ
P8Z1A4Rc8F8PxMZEh93hgPIjz9+y0wjtl+UNUKjxO4MQIeoXxKhS1lNGSAxzwciV9Zd7/OzRri/j
czTspg3MZVbTa7k7eqoxEhjvqGs+XZwxBgXv3q7r1MxfGATOCJAkdldipmbtOeYhC/iWSjTZhRYk
Ksrt9BKXAQzMIv3HPGJCvWqeCswsNKLS6h5LafUiiBvhA/tFzboCHQxaSCCw7LJ1TZqbCSP7+rSl
ysZH3vCgO+Q9HvfiesxEQxNv32+yjcylc0U21ikFp2obKnMxJQh+w4WEy5PSVLK2zYi0EvPPCxCN
JxAcpWndynvY9BUBhJ9bKap3bv2n6lDBkyx4PEjSPUhP7TYLWzri/UfXUaKD7r+vI1sMpoYGLVhN
15XdQhoftI8hGLtE/A4nmWvd0uvq8iOvtiXjuePK7e/ZdLGaFtCumVAbr+lIi4kepkWhr47C0sge
MeDmJ+DLzuVBYMsCTFZmIM3MikKie3yVTNra7lVGEwTDLT+HQtGjiWS15XoqmGaF1T0A48Qqzi4c
k8K93O7zgowJsbBXcDJaX3U9JKzJYCXcCPjcU7PJqdTqdxjl26DhCnWZXyEXIgF5hecIJflU979d
+4OjCYR3R8kJJ/P4kCwZor80xe65jK5JUX3NaqJucreV9IJF9qKp2lsWsCw5sh8fiGY2VvdnGc8M
rm4AXCJ3poCbToPKpJyNyq2xyAj4B6p0+utLG4qjwXLk1hanV8FwWyRzokwX2wuSxbiqN447sedp
FQlSo5e6fPCpaCOaEfLh5vQGoX8nKRmtCQ01DulBhOeWlDfLraTsVCb1kFslsHXKnOOM86or7FFL
ubZ/nRoPmaHEzgBYzAqvxTzCJNnWcmfA4Fk9GI99u9/FbBgHZX8lHXccWm5/1R+/B5dJ1hEJAxZM
benTIWaUE9eetUYi/yZtG2Z9utIu4GF1lWbpnOHqmchQcNSFR9pcShyJjpRIi49m5nRtNlF159Uw
y41mi5VkdG0lWjxLlC2eaNPy8rzcVH+IdJJRBWh+y8/xwe2tyJ0cc0vXSj9EQMXvqQT4gA6M5m/U
u5evmM4G+diwIFQZhd/05lbdMBTpf1bhFDlLSdMbMeFkHd1n+Pxm55Mcz+ajuZl5KvV9BaAHHVFR
jhw8rbKBHzRXzEjeKPxsmo8y42qhb4WI6NSkbGeqElGuwxl0h7E3OUWFjSNCltrP3KShUd4msAjQ
ULdq1J5LMwCyXQGJzbK1R0UFNHWsChO6YoRSJJ8yoEfDriEJNN5vK1QKjkoadVgI5rYhU4BXBZqA
imZz6wqAzmcWLzGFxPsvTjBgQEE+Aj8X8gzFF21L0D7PMz8fJ/HAiexYzqRD0QZbVFIM5tEnIRMT
o4KnmX9VzMTcNTkBwf0GiRQCMkAGlj8KP1O1ihc52PJwbcF8PXjWOKaH1xZ0apviwqXJZVrgIlMV
9mvVU79ImY4IA7UZIhQs79SS4y/PmDpYTWJUZ4LKN/8lbiooojHC12mqXfIQaJks4r14d/Adp4Ya
ui2ZNF5FX/DoADou65KqElHB4ochB+x3F4+7iq650tPAfhPB6XiAmGU3/W1XTG3UomfgyTFpv4Up
2IwgRAuM6AT3p+P27HcokYjrSBXH4GRquvIKCEIuhAIdmXWYI2lRlHKwcxUrIswp2QIhoTJSf7JZ
aeZJL63s8Di0HJge4dmXU+zDPYUku7mZceZTbB8DwGrXoAPyyA4qi19JTeqsHf/ZB2CQNRwhGFW4
VLkdZPVnanPmS2CMYa2AJLiEYZqPYnWx4w4TXGRxcPuwn0/eAzJ/0kvXc8YE/peEf1maAHJuWZwP
tfKd8m1nAdyg4ZZN8qe135n8xAqkvOn9cRNcHLYwwRsYnQqR/7aSS7zM9Cx12VlKiEiK+GmUSVMI
5izqar7rabtcOC3G5cm5Hyo8n9jAAoHovkwuQEjs5OQUiizsfeXX90QyI5C2j7yXBXKBUxrK/Sbk
M14i/DN6vgn2yZhfnq2/1Niw4gbj/2MQkDqRLis6xQlcVKwxP8jYnZB167CMQZWX3JIuMSZLb0/J
wPB3eUlJswXnv9csJcJ+l+t4Oewrt4427TTR3oQEveQzQ2QIewvyj+G/56atyXnqJdt+jXVWA0bS
jw89Si9iJLZwic+XbESG9orN2jM2ubCx0hN6WfcFyGCqyexD+dGmCsVJ5FWAFtDVT1wp7DbkllfZ
9+J96hOm6eF/A3VYFLMCD8zBuv2RM6rXYxwtEQod0CGnITuuXgFnw+21NtLqytWcS6ZlwnKiX7E8
S0hPxWKoqtuJ61m5zH6Y/d8aXoMLt/SuiLHnlFkrH2fBNRSshMPKwnz96et82COrzDPiGNs9gZyt
mYc1uN2PdNiBiKxOu9zyE/6jKM143goMSwslYxd6SNN4wiohqyzypkxizsXCs27vH1RCDKaBqDKs
a/FipORoMXWOCJ7YFKvTkqlpN+NrxM4T40YqpQ2zdSM44jpwYdkNkD0sKtt1N1c++coYblavU/MF
AadBSqHQA7vEsKjb2H4cXEsptckh54kWnOIBbc9v/RoJ9ZBAqMEKqzp7PAdxwh/dIkjGeL3ZQjX5
rFF6oKIje3ELofflp89vpvct9twpOnbPyqlGkEt61uh9JXr33zK7zhkuhJzs+WSKvGuEVrVhTTYX
DamiJkEQem3o2mjJMwxY0IZwA4gFOaMmsB/yIHzGvlVtVzGtEwj92h/kNFo8oLwgQ5o1epsRVL5w
sau5f1/xY7xLk+V1uPO4WISQpWZB2SFfHmk0MtXmvN3TT5wQ+vHXBu7xV1VsEWqca7E/7KSIGRjH
nGYHELbRR1Jte3g7NovlnPTBXCm7ucZOzUTqkoW8CiUbMGFL2Py/qAU2r73Z0Dc7yUkQ2ifgkgis
ZF4ZsAk2ExmAMXLNS5j16tp218ER5wSiTfOw16iK/J4a7ILFWzuq9lUJqBhOgvTL9ipMmOQzwyZ7
La8npA30br0cz4p44o/CyL64X5NO/t1N9Nhsx+QpN2Fm+2h0pNgHlcAHtxesTnV3yAdsVS5K6T9M
UP6yCb+YCF/qWiyNhR1ClvsejNafPsKumpIR/N4fvMyc44rpg4gxu0nCvLxVBMH74cyf3TD7+z8r
/g9E6meKFOyePyuO5RzLneCoP5ZUbBnNODfhSobRKwwvBDj0w2l5kPbBBUrwKYTKodswXEk8kDU0
X4xDyu8DE54jv3LeMcuC1P5x2Vg2aVzsKdVmckWq9fW5VEn9kAl77AnWj9NGCOU5EsfDnN6TCx7u
rmPKKGqD8491hPisboVPIcagU/q+tXJYdM5d8j60QUgAsBxNuQmaYVhsu47JYO6LuRrZpBqcqdDs
Vwmh/qIf9fD49tpiQ/2ztwEP6COo13SQhEczvYQiRtGujDjGn2gstvppLKnA3Ua1IoJTrLw/UwnD
jVO3m+Hyqv1pcd5Dtptw7IqRSwjRHXa+0sr5xIMBtnSsxABWumuaGJkLZwX+YI+51KCaI0UNyat9
kft+ErE2IL4j+KVFLKUJPAD56MivKkMG1r0tgusRwsFw7KiXcmxDFksTCFGR0fA/hgt01TTQb8im
c5KB+vU7W7YvLjG4fTuqM20sTq7WFShparKNnd04a313qUKJi/42khPOR2cCBSGRegeGzL97ztsL
BJhtTUhzyiBspwLGws9lACceRMCrbIbT9qgKmGDisXRhVa+8V/xE829RBaciDgZPtuu/MmOP6Y5P
PpwWYZ6epPCyOt7HLbP6i7LjY0WLDau4L5DiX6gQ7z8DM6C1vP6NE++RLROCc6pH8gghJ8+54BV7
ZiGl7PqZAFz8VfkvW9SO4e9yQ2quVWuuIgG+nbqajSEW3GmWl1yGeHbTriyvwVDrBp09qK+R6I7T
kJHtiKkbPmxD7ARjzzBEit8mEPLs2Vg51pwMnUSc7Iu9FTe+6iov2vNBlgiDFhlGOePWjGjUwjHn
Wr/yE9icPkfB5fSkGtq/BxHge6bl1m6nBvAE+hJ4IjB56cc5K3axfEmoePm7lGxWa99bD0rS1H98
DgxapYjJVD0cgKbF2TcIclpXLlYqrNlrLO7HxLa0fjXwKNdZ2atEeyODVz5/QZ7+C0nI8XVQ7zWt
B70ARyjZByA9CgtDm1qmElh6c592Wwg+Ai6PVKmtsbYUUIMnSAA/CxyB76C8UwmfFeAaOZCToUW5
Dk+zu5Hgswy0X6+SLaJ05S25yEtbJcZYomtG4+yVxQ+c1oOmHbFkaOhF5kAEel82MrK9+uJsqMRB
uURu3YjbJghnXfd5uOY5BuDLruDHjcrsbLsP8NZ0b7gRv9nRtbSQxEl2RL6a5acSlHDfJcxnOxNJ
zgzy/fB4y519zpM7R/5SaK1SvT1tVhe+gFxxx43ptFZ+ikqMMJwYPQekyE7BGtZ72uJ9O+9lXGkV
0rOXwJU0oSmDAJ0Dh7Fc3rWk+5hZ+GdlYoMnptZ1ribEI+HPcRsqGec0IWjoQkxG+4p58EBEEYoT
NoIteI/eqKdzaQamIS95if1hRJaTYp00DuXpItv0jjEY1GBZeR2cTlELgulo799UNl7c5znzazdQ
SKBHzAAl/NLk7yRvJZUtW10+1C63l7jsr4O3u4p0DdTwHHkVqam3eHt34SdJcZiU9X6X1dMHBrMm
7riT4hvcudhtBTD+FbBhlhFfhVJ6DGr4EirqS1nxxXeNIaAIk/IMwYLyo/tWwLXhPAJaIux2ylpP
s3LjqHzkPMNc5zcvUH8kIfM5Ml3N/dCv1LQuaJSHqrL9arJTEZ7AstW7ye9JW1WezI8loLsFnlML
YZjQJEzzJF65k2gwTUJOf7HijktBIgb3+ZDF3KpDqr+OwMTjwWpGTbqE+ulxJ604YxUwb31IUnTv
DAyQB8SevbJJhCm3DvFkAwchKT8yInUKubVPPravepGKwRHyrEF4eotSmc74dn6N6rmjvXqJAZdL
wDVj4ztpyS3/kNXi5Tw8s82LxZHucpFPW7e9j0DqUrbhITZFvR+/t9vw418UM4vpIshLGN/1jdqT
a5ltD6Q7nxfWlgw1VDJJzTqNEA4AI5Hvxxj4MdQRjvLCxInrHsqgTJCtL6qyOj/5GBdmbfKjod7L
stEX4iVW60tA5+VGMHOrsnHjbsLvQEfQ81BDcMKwSNnW8aWJIkGSvz2eu5g0ZzNalErx02a5Uxbd
9CBPVkMVvvhLtehZMmNTv1fLMK/zQAnLyN9FBTfpeKpYk012vsUB+mP7n2Uq2xznYGWVonx/u3SL
qPsEld8kgKBEFAK2bn6Cnw/Zy/mqZhWn/it51UzzaSVLaU6oHRDG8IXxgJGIPEvBkMLAN4fCu4HD
fvQCwD4XkrXbcJM0Z2JlWgT9PCMu0NkCBWi4lD8o964DTTNLe2YLHEMKYHWOaVxrbbaRiQSssjOd
gvzDHrqCAGP77rW5wcyQB45u6YWvQVLeLiwkSHFtP4aMGmuUh1qwkEPR5hjqgdtT4hw8eeDk59p3
S9HYcRxNbPRSMpYbq+g9LkhTwTBjozC80MqaviMhQeE67/frzMjINihjZFXpXfmd6ZBHVdJ4oqUC
e8d8Dvv4PoipQsp5Ohd9eUemu1ugF6v1RxOfiL66W3TbL8fz0d/bToO3e1A1K/pP6JuQXOjFSbWC
if6JgIdC7P8uJopbfiNILlpAlKMQNZy0jb7yc8CA1F6VvdxUSgi7rcNAPag2j+VzbdnWYVQorxrI
GCsYC70xURdUVqD0hH7UtaAsXnqK+NO3ajuaBuD/y1CP7OV/VR/FUO+vAtBHUDQXkxrb7AJFB1Yk
nUHJFcYUCvnpEB6v7i3WvJLXgZYJsOZHLhW9qugjcf8WILaNjG4t/vCtjSji878hFmSypmx0v7hS
Vo9p3i2MEQOAlsK939JNdDBESeAEp51LfZzk+uSJ7PEVfkfp5Ac9MUtC3deWBGstM+14GrySus6+
6IE8xvVFJj2N1ZGZ4RwDJcf0s4M00yrD7ZMJ6nNUOBv6WwztRFhnIJHCSBC+7dWOLCtpzrqO+oOC
vGRyoHdaVZvlY5VoG30tNbY6LzpixUuZ2hsx7VzvDV+DrGkr3BGVyTSnYbx7b/WvShugKZI0khZS
Qb87z0zyPx9a1T3x+Me+soHiyPugFtis4rGosBzXq/krJl2/FQuvZupuSzXIDgl0248KCMGPcUMh
IcXc83/haCe0rsfYuSPXXEmZP4YRTotTJuFmbFm26TSa/5LPQGnybfmaC2EZsj5D0eMolS06PgH3
DsJTRLd+1XHME1HEK1a3PkA9Wy6hguMWLZScbRjDu2j18JS8WpkARsrSzjd+2OxhbYZlkOywMWPy
kfFwqtX96Be+SF47C7eLtF5ajb4sqqfS9s8X4ZlBkvNDse2bgokyHdno3LnamU2F1yI1REEGT3Bg
L+m2Mgtau35OJAA6ShAWR5n4MGV4TXCnbfsLd+Qjm3U0wi7WTzTTWeZL9ypX6TpYmTR8ZmHKk9Hd
HK7VH0biKFAEjSlBevpMEBHoX6zKMXI8CyLNcYzoLkWkzxZMgMkGAyvZO1eEaPlHt62fifmSH3Qd
Z2kkoO+4r4ypnl8KSFOVu4oxEatjwyezx5hzMF8Sblo03uccfxAe60NqA6+EO5HtiodDf5Bk/pSx
ntV3sk9yJq0JSnfj/j61XKh8QJO4A6kUZe2YeQBY7OmlPTHdHv/pDSNBJvEw2GrVXoZCayILXaui
MLgT9aMALPJO6C4KbTSXhlCZIwh6CMX1KotKeiXd3rBuf33ECwiG6B+qnmlwRzIIv4RpxjROB5Jm
7NTD3T8v5qyAtD8NKx39ZSSeqaBLY4xhutgexB/1dKeuq3rJ/hY7R15vi4r0QfeNmEzaCVugr3KU
LWBWXLagBcEvrrgHjYbYqR1VU8nJYrUV5XgxAK1DUsfBHa+IK8VLl3Xa4vR6Q8Wgi9uBkTum98f4
V/XH8gVGK6V9GCev8c07+QCd17BoiOqfls7agaYNIUHzYFkb4zhudMEDGmav7OxM/KmWltwD1Fof
poPMsEhYXP8pA2NpJPsklFZAGJKTaYRgq3vWhF34re/Q13mrtTj600w/Y3aZyteLwgbEinW29Dt4
owMFYinGON9GV2nZ2XZch4I/B3N4YiNhvx64LJmZiT80am6XypQYkTlqwSoxAYQzzDeCxLuYYG1U
i1t147JGaW63eehIh2mr6kSGwQ0WH2tDXGIhYESiLqtgd0SFsgbh2brOl6szwkvFk5hHMkbwcD66
0uqWcRll2OeQejK5j0iqvkqHVr1Ej/m7S+1SU6je6PCVq5EQBDKc7236H7ZaUde3y4l+zByN99eN
mznOHSigQ8gPfy9dIvGTEc1H7oF1aTmn6VvSLAp+acL0jfZ3PG13DMSiWon2Z6u46Y1eJbtJrWV2
+O2u1yC/qjNpkTifG5j41wXs+DD705NtQXznjLgq3kmcaNQnVlOolwZTb1B0odpTBczYPiNHSYoh
0il2h1aSaCh1Jk0T2XUPuB4nFWkovB3NuW2GZNTW554m+pNF6HvIobJ3iQGvGnKyQDMO+Wd0w6YQ
zNapVT0De3NhvPHVJ8Do87seie0b/nmDbikrQQZXebcv1t9JcuUP1FWMcelHFjTwHl+9jncj0yzs
PYl8Sh1P0Ry6BApsiblj4iyhAyzj5OE3IabohagPT4DkQz4a5do6c9fVuhDPot2US4I8I0O+fJHv
3pNk6bM3MVLC2Ip/nJwHobxvsYW1axr2O3PxKZF9eHKRet9OyyPjtyJx7vqjsY0X/3vmuxEMlyoU
N2lTsRfWiLuGcuY+AhaMqLFGs9iYLVkljJeIGx7akvNZ/pWZGxjY+bjqvUfe4NC2EplIDbBmNlvH
v8nQiMtdfEmgxq0ULRJpk7ay64fGEYKPANMHYmIyDoAWnBuRBg2R0pS1MM9PYRD62W7HF32bNv7S
/2q2D/FpbGEPkePeh3rKEwuAEV0Xc6kKvpt9p2BS0t6IgMAhwmahM/0equf+0MkSrNTTJdxznavr
cW6UFMSBk1xwS3Lodz69qEkyRVRQCxWD/WfEKuTKqVZEZp2Pyd/ymXCmrWz+kKXqSP3onoc4SNWY
TtGcWzake7AfhqnSd7DNaGTvd9xmyxEGozmtHIgXxfRGYZW5CGyPeOPodPCjZTk4XTjyh32EWwdG
7zrjsGbXVB9g3Jee8/QsMTJXuSkM+xuco3HMBETygZWzKl/F3ZkG0swypjIj03Zro5mATSsN7+E0
VB6Tmk4a8c5LvyW3lMI+gWb1Al/X50PuzuzTfyXDPpX7rg7t9WPz3rjGQzZGwTRp1tvfDrrVlWBF
R8d9mrCGdZBnR7884uzE2LMeaxz8R2olVuQyFsK2EeflEkTGUWDqn/yBcuxwoGLQ3GgmiKql7FE+
ztsPrYtWESdmg5Ib4CdZ2fUAXB6VpxkacY9cF8EXHL0YkvNRc5vUNlWSf38bCvqIyw/rtXwna1Iu
OehDRkPXA3QD7ceSMoQClAyZaar2oiCozVQE7WRqg5VZ+lzZP10EBdxuXyHmpSIPfJb6VOfrO7gF
BhnJTtz3NJqZISDfFAY9aNf51N6opiRVRrKXMQu3v7FP/Jkv5aUfcwZ4a3SuFfnrqhI6RKlqCfvE
CazJ7Su4ovzbCtUXGQRXzBV3H6K8l06jbHDO+ftDDCBAAMRlYZIJwjNR4MLVdeH0dWp1awovDBbG
9faGseipM95aFhxVVkFUhnt0wwXnHD404zSudehSsWj6mYK8rxDYpIPbL86c4FzlrJr+PqkQyW2s
3vMKcLzWWarVbJX0NGfGZEHIRNzaQgxq7sZvlTmfuu0PJorw8vv9ZIx1qgezP00wmq+Y3NV+65qA
QEl7SI0mSixlyeKyFJyJGqkQOa977457Q1nWBPUCOQxFhP0A6g6hB2LhpRQuBsprhRGwozdtj8jc
Xe3e5oXIAvbrfgxzt8xOiYKTN510pQFWGD6VM9DO9GEX0XX0mkfwrqPALe1UBJ59OByDOF+Rb7md
dh0xFL1V9m02bV4GRPqfs0qVExL6FSAu5xeHFW3bYq0+KintY+5/61/TekiQrB4xprExz7pz7Dso
rZ5iVFappgt5Tf/TVdbF4N58UJSrqLfS5YvfN3T7m12y3td8iI2MqA6vBZezebmkpftYUsBSCuZs
IRvU10cDtfl1VsHMRVpbl13ccEN1ilNQY3sfRD5lKstRyJWT/8mNc6d4xHeBJWOc8b/O7GJMGA9V
03JZvVEyBFukUP7+bP2ktNCHb75z4FaUYTE1JCGQuiQLjKH8hwvBa2OFdOdZLXkKPBADFdZUkNXt
xeDSTXmx5GNHC3ucKPchaPGu13Mk5bf0kBKD/sdokV3iVoESyQILJSMvAuasXD2ymuodHOirMQ4a
HxK18dtazoDVYzcolsz0PVzsx6gX3iIdYS9HW28mpcoCKNnBkijsEOY+UemsRQTRKQloLbMCKKVt
Lu7i/L9VXkf+8Vdhlr3SjGKUvb3EU4G5/jF8g0LimcbMM2XiWiNXi/Z8/C+SyHTEA9iCBfyq5/qK
VtDaRHS0qiSKgOpCH8vY1MXyvfnumHIjtMY8gzkDwbgdDJYeSucOjxAPtZ2GhrHXZqNPMmVEwn63
lhaDfhr4Vz0yi1D87ivULf68+Dhr1ZK3zarxtW8xwzb0J5yvtfjUeQCM1X5BlznJ3JWh4Zx/m8tk
zfDR+n/XBNfKTuckZl9hIdFLlr+Ye25gUUHGvf/K/SvYKRsL8Psh78CVJ0ai+g1uQWCOg5kcF5qh
pmtacQNf/n+T5UV+b+130UT8RDEPulsQ1TYgl5Sqh4LJXFCB3wBwKc+u9mLo1Pmn5apKBiM1nGm3
vaKr/eq3GpWLKEHoFtYCgp9lDE2MwBBqaX1HDAyL1hv86nmn+QNaRrieNomAp7MHff48KVSUKeJI
NS51iNt49nMX3y2jrajWnnflAPlRDr1BwWnCWjOMfUXeisbY94Pi/AZ1gXeBpq5FXzZqdX6K+MwJ
z6UdBXExpUvmHxMqQRfPG/CXI2d7NpyioHacmNczkYKCqKt75iGYYczJbgloQ1MauqPvY4qPsi51
ViMPys3ADreuxPg04jS3m2ahiQSHlGgdTepGShKoCLzFAmAhtGrsRcMG50aLEDWq9g4g6wBS203g
GdE0saPoKN6EJK2Nl+efyHNwx7T8sQIpmQA9ha64MZsgorxEYZgI74LQd3tOjGVd+Cx5+MwJTPnb
3E/fSckzyyb+064L4Hn0wV+iN9XMXRDjvFY8loF5fpisFCbTscAsmfjHeF6vkdzycF5inaZt/qT3
R1AVxSDYGWSfdUg3jj7pZqo9lRd4/QSYnqCVNPwYPCGVNy7t1EXmz9Dri+J2L99PFaarfLnRtAgm
tVg/NpQvv48els2TfRSzNfAf/AtGBsJCt9TARZQC6LrkvxD/0/kluNy+R92Xoy7kPlrdRn6v8e6U
2ahHgH+CF4QOkSTpTLkPaVP03bD7t2JZr8daMlHt9YyXE9ew6iHfRgz6Y/fuIuQIeHnYsotgwNZG
qBihnEV/yN7B9SVKO4gKNaMyVv5b1P9V1aL7VuvkNOgU7ZhCcNJ2fwXaXrmPAMYZOaWmqFOPFb44
DK3PjmarxfKlF4we9/7VKgMkI0x94vAup31RFLmSiIpkYT6VqQR3aRsLfNNKMGmw2ZZHd4qFQjKk
dCrSmRPPOOj7i0hK7UNPhpgY4+wNrdqRbhLV1DMk1lQ01nPGOldw4crTjOvwzno6HCHEX2zgofsx
Bhg3CORl8i4s9jxyxN+TBX5xHvgUeNxf3/DiYgT8K6Ontt7frDaJu72OwKTvlkYrbGq0Zm95/uOh
WgLDzXeTkG08vsp/SRYfhnt0KO6HOgaYDsekmdYu6HeC0BU4iLACqAW4Msu2C1c6zS9ncDhAJ1Rg
o7rg8VGEhdwanloutySX4HsdfvF1OU/0skDphoRy+7cDdtsQVjHv1X5t2/ITQ//IzKDt+FVIjSR9
GiXv1oiJjpLz0C/WJXQbojDXEnL+pteOM380/A6h9pg3i1cC5twULPvRQqMeaoHu9u7Ld8NCgo/r
prw88NcFnTYWRFI/LQ2vwH2cQeJpLtQVC4TILzvQZqdVyRDdXYjVBrEuP+P22P+FZ4Pq9rXMeZit
jG3qyOlLE1QdaAXAT9cxTV7mCOlK556/Llq+I2s2taXfqpg97FwK6FD61yohX9K98tXTAv1mFI1Z
qOQsZwGJCU4tQmMNdBfPG6WJ6fp+kCY/9MMoGFBgA0pPZiFm9lUam5r7YxJS9I9RfwfwisWMGMKF
kEKjqLaHmraXhkNG0P8IKPOBjegLZTDQ6hlmIsztTRBQRr93GpCT3FRZ3Qk6EgDATXQpchk7EQHX
0oAMglXSxwoJe+kGlMJKBWpmSBP8P6KYv2w6D7hbKjkwCYSMAE/XaW8Ps6jtA/N5FRw5F2IL6q+A
39aVmJpl2KfwgZReNQcVAfziIN8K3ozxFD+iDo4kzn5+x/KS8MrYQ7CWoGnEBh9WUysH2ya4ZYXV
uxM753iQ0t5CbOVhc/KIOSWweNjxZLnIy9VX9mIK+VSN18j1i5vmAh9JznTjAHJpdSjmXQtqHb8B
WZdkRcteP3fJasENw79B7p8mOZfQqljM0FKJLofy30iYRFxVWQcgPABE5rbdBifsCy28dYKuPqaC
T0CKaYCPJmNk/Pvp9AnHyv5Xb1EnblVHRk2RMhytuiqwfbDsp90IwVW+NyGlxuu9rN5jjhfwDu9y
rKBS0oFaL6tcZYbUUtuAgY6kbc0pWK7HHBjR0sFodKFQjgB7Q5+3HfdrmbsG52GHocnywQJmZPHx
Lcqc3SzSho6T33IocowQrKdmS2cDuQTA26b6UbfKiKVrnNVuHFSpAOrOAGtFuNB8Y1iJO6k7mLmw
kztGukfqR2Ofq8xSSIpUo9bZ5lT2AxMJj+mY8Fj1lkkWxG7SZevCihbVxWtNUziJ6sFTZBpD3fOC
9DFK1WMeBhbCMkva0qT695nKbploMKAp/JGnGAEtHl8y5ngldU0IV7bjMEWj7MiEfAbwt0YVm9FS
UEPyxo7vO7oheATqf0eo88g9dx4Qzhu3fNVjLjd1Q5RX3UzUZM3p4HkDbnVRzCwoxRSH905z1/ZK
TM1yITs0k1elM2+MnSPn9dA7a9VH6XRqI7GYnvErxeouWl1usmb4NX91tS9wtRduB+j9VRZQvUcX
TZoK9IZPLV76Wk6Y8VEFzTIWSilkT2JIrtjHRfbiz31Qg0siQ+iTwbrfVo4TX5pqDX2+63t+6PAT
FYjQK0oU0it59OklgEvwW5OCa28ik3Vyh7GgGED9Sihd3LQGpeKFVTyALQxKUTu/iNeeRuHOt4QD
ShM9cVp2tnwpTbhMg461SsEpDPreJYMI8TL6f1o5pRNLSievwDUuHtljk0V19KtY3MNq2oB+2mb7
3SDmifzkT1nMtvjz8VaKwceomdwELtZMvkLphJqrBKVHVVhfWjMBm8mXYYbiyjkUJq2RE6NWczIl
LFdAYPZ6FAlwPFhSKdcE+LyYtduiuUuVH8ztNrTNcmIU3v1SUTthz8lOzWitpj9jx+XluylQsCPw
DLtCqnhCsTu92oUDODKohUqUZYurWhtC0ydfNYcoF5U/zKDXGyHNMZXd9kBVhDQ8LMejIbkSBivw
77xULJFP2W381O4bQqB0vNININsbfDN7Uzk3cyCsggfl7aGodoYm1U6GnGiyC9a2Njb+3X/XvKRI
ljLPObFn4uckR7bFqguRwTjc8H1DeWu3TsgkGVG3eOzV9UnMvFzj2idFT/MLiv4+ULiIEKfqLVm8
34epDy9qmYl5V+0Nh7BAG1nucJBMj/QpXIWrTAE378e2YLpDEpkKAs8B++iLwUN2Iwrv/D9zB8oz
QCjEaCj7Db5DYJ+HVUezfPZmu60Sl8z8ok2lhXoJp9buae+kpI1ge3X9U9hRGUoPFplwZVoyX09H
C+XcM4aEYDnWQ0FMhSk8R2RcqyfR31C15e/3C5mMMIXmwRtKgfsv3a8Aw7XCzCWEVM92FN1H1VoS
LFaHmGOT/iiVupRR20ai1t2QITQEgEm4GWfXEr1CPIX0DF4dVOJjt+Lyrx6VP3sjhlF2GusEyN79
w7a+Wp9vzYjSx8fc+L6KQ/yWKrA0uuWA9mQT9HzMAiJ/lAolOUzhYD/wO8uJ+XJwn3R9CYtIUdRM
GQyJUT5FPkpH+w1R4QNC/AXyPsEBmPemCARODEWXmarrg4jwihUVj0RBZe6JlYbKUk3Tw6loxYQb
VtKvLxFA67AE+1JBK05FdQoCtrQB+5ZNVLur3YR7c+XjKcvQzSwq+l2Yc6CNeDGywsWm245SEZNn
ADQfBvB2vqJ0ItTuJ9l3vogfVdZoVdaGMwm5benf680CxSvUR3YCa9PsDO28j04uKekiQ9Yo5qsO
qDA47bF/Oi1UZwF5bIqZ6wvHp8BRaG8Kv1JyPBWwhFoTCfPnG+IhBvKDTliKDzAYUax7N/RSZiu4
/nrXRVtZvD2ggQwk38afSPfX6JmVTPUoBnu1QQdKfH4P1z0wAtsALixN2L1SyaGSUUz/eLSYEtns
C/Lr/TvIm6dvJCkk55ZGLTVEJtvhPGG0gE/PeD2PQRHTdM7NEeAVbyg9JG8Kuu1abQIcixSaNUPn
ggmgRlOe3GwltwmSWvC2+N+TgNrm19mYA244T8zgVMZEhfv1xLP+7Oz9J6r4HFLh24XWp76JrHgk
qLMg6O/GlGcaoiFvifRui8QVREGwIwt+ll3WM67P4PC6dWJkrzMHXgDAD6+GEEsC8kNIt8HKQJzf
KojXeb5NdUMo0YD/13KT2hpjC+z9WS5ISAFjW3STCLR6BeKBWE2dbu7TQvV64OuH5rsAN7bVaDQ1
ebT9+6to4ZXsTJr86G/zN32rmwTMDV0F10PyIYOEtM9TLxl9a5kdlc/XsevB5H1acuDLsNHwdkCc
UdiuusWCwiwwvtN+JAs22pghoWPeQAeWaRiyvvKtPdBeGctnGA5EA1EkrOaC9yTX0EW7tLHdkQXw
okitiEODKfeWhhWBDxRnT99I28RdkAHn9ZrnkQjBSKoQeBSL4tbe8wRe5XFtsEPuEllUp4Q+uUYZ
qUCICRuzHZTj0dIE8lN+uDSnXb5llw0o3l/il46lOyhYleACsPlrisrIPacQaYrSt5NuKSUisQk5
IdAYk3oveDqbi8NMpwZKwDC5oCmwvMwL2ooUmzqeIL3de2n0wOImN1LNp67ZbFC2Fw05gpl6bWrM
SdoX3JKHnFBckJ9JLU06bmUjIYE++WaFiBYTdbGAKwSiwnzMTI4gJSCctPcnmy0QfI+ZfGh2lV4z
SAYmTqbI1y67bTYbMbpWMHWfyTxlY8smXuLW+d5nnTIvffNTZgynP7Isy+UMXq0zRPorLZ+AYqHQ
CwVAs4TEJOnXVvPnI6ITqcpnJ8LoOrvb8khFcaxlkMO5YhxJdxoBHUNVds0NxgBSvb6dGQzYiL4g
PONCdRdgO+4R3YWFjf9o+jBdJsgyk2zAmsr1qI0qIdKekt+gBtLZYTURQMGzUviVlqHRwDi3C5J/
ykqVR2nzd/kw9UPM42H7MkFAotquQ5hq8E5tppsXr7ZdiUWk4QrhgOHJ/YQ725FlNXzMNuMdYGYh
teQrDxBG4pPaA4FoOweNZTXekm2sGctSilZoSbGTB9UAwc8W+mcsxVZP5dQxCjUAHeq83QoU8fpl
UXpN05p9wayEQ4M7TIM8zVsflZECFcYejIPM2DiDX3a6zAK28slWKeJl4f+cu1k8bUM9HHAIcHiK
qPOxq8rZpCPkFSnBAqZYma8bJTNkmusY/mhosQwGqff7jbbVtLm5UIYdvyXtUMifoimXc984yG7i
Fey4zAteO419DMj6vnPx09U65l89MqwUyCoSbyL4vev48KUgR7d3trkDcSH1WS+QSPzLS1rwb4cm
WB3EojtFT8I+epD0dHqJsfl6socWKM0VYmW48R2f8zcCie7LBoFzJTom3SALlTCt/njPhawYALf8
XqrvdI0xCFkEqmkXg/67TE5sqllLihGk6Aps0MhHE5nBJ45frbnDeyJ7A0CmxpVoR3JdusWhrSku
PKLJyjgD46ufQhaHv0Nl/xOcwdLtcy9vhXcniMGvlJpbmZbyij/5NVqgNKUWeNYiWY7Ed3ErDsR1
vDj+SGl7WNMHbsMxS9I9gJINne1nxLsgZZ5L6ktuxKz1veQZZX3JVXyLe4+RUYaLDnfBPSJ5f4Zh
mN8oyZi20OXpgU1tMQZj35MUTpaOC80S9LgPnNZ4mOlO12peIf7CzUZ61XHwokENBMNh4VWCONiY
/h5JngkjnFeH8Fth6qvzW/VuMMoIRsb4eE5qHi66c/LVCl2qq2TI2QplzFAu3TZij9exaW1cCf+1
cyq74tN0OO+CzRFq0bByEjOPK4OymszruCsDORhZjVvYJ6DS35ai4QFiPKoJeJKDD7sLCzI+qwVB
a6cmOj17Qe2WgnS5WyaMxfV/+6+MUYlrr1ZQVtqtZOkBNz0B113yJhhgi8Ll1aDcV1pylWwIOkJm
Fu79TAv2UW73fxu++tEbhBdIZ36oI3FBR0fVSmhnESoVA7r1Ry5+fBci98SgUJxTq3gEPVRP5oea
UYULUMycXeUj1Sd2gKZ/Dic+IMlPn0itzGy+nDFy11mxwQJTC0j3egeWCGF0nFbrKifl0zwTzwFj
WzvdAnCVOqZl0ERFycmK046515yaRLgOrHo8DwLbtHGdADvMiJECptWUlJWSumkrVyxy4JlC+rU9
ma62WYBu0ARP76dpid0Slh3rPA+x1okqx7tdpNLACvM43QeUQYv4KDq5QNXVEs40pxtMC2HYbB0U
VN9VB8dFJP7M3LbsFIFMPdDuRsJZGIBOZLHfZoPaWoXmm7CQhMLt6WgHxEHr56BYDpo420AVBXYo
utxjozx4bvD+wJTUFZ187GvngGEweFYb2A01haiBGvOU+P65eqMk5oViDfFhwzuwsO0uYh3jv9h2
7IKRlIEAkRF0vb8+7P03cEljrdBGCPRhliuUL/rC4nz5SCztbTMl0G2lzDg9uALFogxIFyMxz3G+
LsIyFDmtgSb/XIiDGDrNEhH8rRDFxsejO/iITxHAD50+QpvPyL0roE7e+Bygh3AaTVEDHB0cpx0h
7SHAS3v3X+dm16riO80KSa2/9jAH8O3urizwQV5nrWCykZ0OlaCfTfhelyu1gw+ptX6LJS4Ulmcx
u5nG37J/WT2tc+aQZ0BJ+SeBj2mcqJtO2sIIjXISmI+/3g1ceRvmcquLAD4Fij8roUnjGj7WlTLY
v/eiO3d10m9RnRraO6izK8lMe5spihKox+WnbbmnZfBqnUynOJIsZTXTYnsJ6mJHoxZVvQXA6qzF
yT7QUGQvl/pApyKCfBigp+SayrcE68y5xcPtaw3gSmQOzDTGzKHLaOo8aSVOY8A1QrDOZy6Lv4Ud
IfPAISXkCBlVTZiiI8Vu6npPSDrjyEOs2gfmppHGnRMG50WyVBH5onj/8BZ6GkiI3TeOOC6fU1qj
MhLzC5SGWKGc72se0D/kjjBCDJXziwb/AGtu8AKSvjVmBO/d/CWeKwUPDgi6Ydp4XTE+825/0Xua
j5bL1+lqCcC6YuouUF2iqSM2J+2p/5e+a173moAB5Vo73YmkLOkmroGbyT8l2gEtC7t3oDaYOHy6
cEZ/WTouLVeBiACBcMj8rLD/D5EBaxMeIMwIzTKh/1JbCs7V+b6gV5QtRttJbrDGqwgT7jVKnKtm
nSCYItWHBxA26zhLweXhAb11YzuNqo2swJa2zRSwQumi2pUMFfcKac62ZqBY+E+Qp2ynQPy7w+5b
dRjisLIHQqo3W6tfxFHFg1VVavegjH+80PuNlivrsS1Mu7oxm9lMcCtn6blIybjJOJ4cqxqRE4wo
gsY7Cb3I0oaOLm5FOXiHH7XS1KXGTK7UizrlPv9skxlO9SHl4Bf+J5ZDeK3E0Ua6tH25W0HT2VNb
sQ8JHCfKjfxAiBHNeh2iuZ1vEb0M9IAo/Qkn0r8WRdbiNsHSuKWyErMEcjp6Ay3nV84tgw4+BMBp
IKalcUOOIyzVIjWr9P1SEAfAyJ3oTcXIvqQrvf55o89eWQGYM0I9nMKFQc+jEVbWNoX900KAnP+1
RTe71/ELThGRTJ00xdr/T0DysjyJ6x6BSR9ZlsDdZtviLeV6HLyIRs/XqYG88FwplBN6Dpji5UXi
3NZb3p8ca0WC2xyvodTzIFD5KEwIxL6HLHXcmxAzel0nZIcjW3aKVSHBsL+XjmjGSNL5Rmv7m1N7
4yvYN3MqqQ8LQyc0/19OpFgxV6oCKZng8ebtGAEnY98tB4LKX/U5n9GDWtzkmvn7JFN+SfUEvCF/
kxoExKkk8xWwSR7Af69WV/rBPmVrL/CorD+3PeT/H+hwjcCj9PIMA07J4pPzcnL4LntnirW1Z1oy
ZI+dZBypeN8LVCMNqbAfr32SZq25sb7/LA1yvJT9g80EYkn2bJ8ZJ6e7gew550Ui7CcZpx6gXW5t
Sid8YmEC42/ZrKYG9X7WhRdzODr4mAS1BF1iX9ClT8Lrm50/g68OAQffPrtOit0tadqctz0N08wd
v8+qKDzx9e9tUeBuEYuvieO3iiWs46XFGhyyldmM8E/Q5q0PRnLM3NHbj6KlSE5l15Uy541KqGMm
5LVeiTQukhZb3KKWuDRWZ3Fr/pzP9B3Zi/bGVSOPyEDKbFm0MpJwq5/lNlrgxVXXewI/WsaLsH/J
zJ+aEH8cOnBuwYSkwuKmCsu5hai7MXpr/m0L6aIpchVwsghBdWnPhp6Z+qV2mWKq4Cen70ir/yLY
smv2PNMD7dWRgf7ADjy1tyTGyY92V9Xm+nmvEEphazwxDK67luxFTDAu0Sn0ByVF6bnA3wb5ctgQ
UHNCo5jkNA5eCWzG81o/9/ItGFlU2gQH+WF7fetjZD5GCWxfS/ABxoBFGrVXBJFhgoUkgZ6K76GK
nzHk+xjzylj0ApWF95FJ9yifxoXjC+3ZEPuqW3IC4hPWvkSlQr/Y6eLRoq2QpAprwoQ6lXHR09m4
AlyohWZuGaYD6nOBeyKDI7H6hH+NYdWr03iCgkgyTJngNeiHKkOR51j+aST6YoDu/HpY/0v5wNef
VvJf6fwZJSRQk5Gy5oNMS11t0A+zbyoYIpIulCCQk8jHApOmKRCEAvyZC8ton9BqGY2jh5TzapQm
FbTDyX30YturG/bESns5UFgVvm0H1Z2EzaVEBMST4omKEyZoluDqDVcH0d2CdpkSPj043P6oix5b
/22PQvysu0+NT3E5H5mrIF2QzZR4DjuLv/MqLkkAbFt9aVCO5J/LMeYnCCxYi5NpG/MNy+0LqFQK
2JMHk5vk47m6nqeKylJ+k3mhlTTfN0+FrwSOkgx4absa6LcOLXUDfqHmUc9os648yMFqp7kosbfV
pkVQH6qcZoLGQqy4bf+greyNGeuQUN3X78Z9I94G3XxFWd0DBdDQiPxXsQl4chfjD7cbYGZZANlI
5tV4BRcaChxPu1JWe4LWOdZCuOGkKzwUtvS9MUyyVOodTfEc6wUwCtMwywZ+0R1bqhxIQlygUegk
S5B8TMpu8DYw5uqgu324AAfuu3EoArrjyoSVcC4yJqHubtXwELHfIX/0xki40GJ/E0Yn/7BpULfS
dJkalviuOtZ1ETLyuXs/TSUpe489ckxftcwwEUaxM94uBBGMFLBbvfVRflennMn914VX1ofGDoo3
+xDnoEn5IlLoDijFBaT5APc7VW5dD+YcntNZG0weD7kx61LP/L/4NrmSNZNIZssRFWZs1h++RGFV
oR8uZWfX2CknlqVIoInUexwT9efrZFNcg7h0fmiYWZsES3cItAg2ifiNTAnrJ64ShEOYL0LcBMbt
6p9Pa+bW7UHr8VcKC2AvmSSHHCXJzMKbCn2FZNdouzEAqHiG7NeT5Z7igSbzcggQuxPjGZsZ5rY1
Iz8cPGlqLuRwkAq0vLN8llP5P6YxTPFC86YQ3LZEwl0EaKFH6hVaumw3gXsGGIF0DjIJm4adYiYp
oyPDRj/+ko0yacIFXuB45xvCRW1P4ka9BLo6YO21qsV8aNrpKWT/Ho3y2WCES8NGYYuH+b6ww57P
RxYCgPStInwNrzhzZL5kMYqxsOAH8N+RMZw8czPaKG8jIOoDK5Mepno+TwbtSXq3BzK8pSr8rtam
4aiQEHr+Z773GJgD5F5Gr1z7cuJjRso6Go2oxU8lzIcxJpiIDRklmlQZIqcXeHUS7uJwG+gMdRWj
8PZEMKLqn6fju8oWHY4vxzdrBoHP/mT8WlwU9IwdyuB+6bzs5VGWR4pC+dnIgpnPl4iC01c9rhjj
eJQueEe2kz3HuoOrNbV/VVRE/E7VNCF9Ml75EQFKqler7AOK1Ct8aFiR3pAY9ROGc+vhC2jJUNyQ
KsvgDjxgIzii/hNb4oJUlIbXv/Rb60789u4o87c6pk3+qzTC+DY7RC7e1iRAFNaY9sXSIEZK6X9y
fM+Z5V3vZixv/YATNU3XB90mpTNRShdgtA8ybQZCaNvCDwJe0BPuusre+u81dNABXcX4hT2Bl55r
XMyoUxpteU22wZFwLljXfFkO8T2Q18AMOOqLhex/HsrBS0DjMzzQ2WmCiqFb0ayRN20o1nlbp6Y6
Bn6zC9lZPFwdk7ILBRcLb2FM003nLdoDbIyPaNxitnQk2YFxH432+RtfOWDe+31wx8hMCei71+H8
DGoOmTCVe7X3SFn1GPejTRmwb0LgNueyM+87gcUZ7tznppyuyqD8rz+KdLXORVcubRer/bsMC1PY
Tn9RSpoGMxUkvga8HT4wOXdGtKafTequhUtO06TCfph4arFI7M6aXJOT2G69/Os0ZqFXf8VH+ugl
/kA897Pq72DNUqvcJZ5Ho2+CMVNGYkTXJYhR01z97EIKfXGVFZ4y6jLiPYTEs4J2cRnguppsFFSr
aPpd94L3mzwoRpeuOaBF9DGVxqu4SGogDQj9HLBGwFDgnUwfjOCkfBHZgO7p9p6stcLw14AxZR93
RpBCpSYb8+5isrxf+fOFlEbw0XUV/E42Oka0v2HKS70srl1iJV3/ATb2gNUPV/KoDYamzvUiD3ye
ciI72tWlBCRY29JMz7CUXjhbpJQQVHGwidNtX5hCOEjv7z70YZuLFNzPaKZ33vFGy2/3YJym/cjA
cLNC/dmkGMKqb6O8FYQHmpnOSyFKbZ/YgGkOMdi3pHNd3MO/Gja+9mn4j/mRoeyzBIWBG0DJpvvU
55tpQtA51LzvUP1YxKuRFkSOpoRekCzA0TaJO7ZVUGCwL8kmUSSOaDffZ0qMKgjVNYy78eaOf/Gh
Pwi5ensa+u3nIrEqsRJr5PFqgnVYEmAW9BB7K/ueyc5FIqZD9fyeh/gb6CEXNUGtZ0caOAFhVrNg
Jj5pOxd8R1p67B5oXHmdifGHlqCUweHZrsrkeNGWBFZZ8unlVOrgOr5BFVfmb54VLmKyA/mhqKSE
+53yhEAN8WPH7aYAqkhrtB0w0O9QA8jAws/syGPq87jMeH4VM8/Y0Zztl1/9akBIBivJldjBxCUp
MmuKPqiHsi6ckG6u7pdecq95MrBYBIax1r/6ZRqpF6bhXDI2pzHwIvi1+KQ0C7mRyJQ/kZBlbx4M
k7EUHTrYbcdftDmXHts1EK/RRXkSLCSklQImQRqXgj1FhICY7F9ynrHaBMxwMkN2Fr5U8ecgX6Hz
WC7klIj4MvIXs8TO78sC1NU7e4YX0ybatszn5dlshr71WeIBQdnSv4ZGfu+TuBht8MqjTJbxdrNk
wpaH0uRl3FuQc3p6O22VhLGs9wH8KCrkNwDXbNTtolfuWQ3+36tXY/ZxnqIE59S3imUpMDO2ImPn
yTh5pLBovTy8YnAsPcBDBLnk7z7LPODDlTISy+spDWYTlwV0g/wgheu0u8BIFBJk/zeK/mnVuUCG
LqQ1+I5gn+RSOO1WBdEknAXhzVR003BYBKY/XTXyBNtq5kSXiTMqOGGXvYhc+ztwEM8r/qxCz9/6
pCTvhB/5RVUvD2Zwv3lOArAAuB6TVE5+YO6c+jD6u8cueiWaO8NyctU0585laaoH1Tu1HsbDiHnU
VsbXKkwNFXfcZfLKwY1HQfRdbWlFo2n+NyRSV11qt993v0V0KfJ70m8LwWcg3CKSgISHCCifN1WT
FZux7IsaRqapfpq7dI62rjZzJZtOhtMZjuGhwOk7C4vsNZY7MWszjsvoBviZ6CyHiCQ0/8OkUBka
JZ23kyvpgaQPy/eMeG8ndhopfO2YLzn48GjVQy5gejA0qX0NXhVewHK+zdjpkS8neNJWW+XIKD8I
RAoRQ4iLMRRDiQwRxnq3EzWuvpji1cUJRFpCB7Fmp1OJz4hZg5uZNzvY39iim4XTs3LHTG1ayo25
mAs6ivWnskHfd6chr4mkiUXJGAQ7OpxJ2SVIv1bNIjPkUKQpsd06SIhiTcNTaGnaffXs74i9oLUl
9jUC1+6E+ULrXHHhzvZy4TyTaoSHpVJ6Zi0RrTQ6cvEoAjbfLxwamRPPsKJC4oTpTh31PS71b+yK
UhElEQBHd03CBjA9b5ZK1Ry3l9Ur+lY639LuUMJQpzha9fXbIHZ+STAId2aD9J2TnqBOt9VbcSqu
CoJO+X7brsXWOkD/P/Ib8m/1FyaHL7VQMTwHIhbipHqLGRg2NQlqBZeqNJJRM4q45jcRJzSJrAYf
b9JC/nXzk20zgc+HtCgmkYTctH/nH8rUu0kojcBgEfwp8FHeelri4fymPsyTyCwyE5udjlT42hN3
p57aYuiqmdWLrIMPhadP+5HhEpZWe8ganRDE5m9yedp4NBSrPwMJGhTt4OVwgWl4H2BG2e1tghJh
heOHnMRY1RenxCg7CdRCoOVO7U3WtxxTsejNZjk9Gg0f9oSfjd/e8+wDv9J+5/0N5mbWj+w/O/y/
e5GYv2k8RfeN8IiBk1pvA91JxO/C0jZCcKgSTP74L++7bOY+zB4oce2FNr0z/ADnDjjk0SSknC5K
d3UTLcOWkcphInZCCT8ukQABx+HSM0wTtRoMHoNe1vh5wcO617CW3n50tXCkYRylV5el3l5flyi1
NC04d+j3O7vdX20nyv4pr7ti3XlkBDX7aJg5+OddRK2fmZENeERAmIaAxuDsya1vQEZpkQNVVKIa
c6JeVRVCX7P0Hxv0LVEj0CPP6dftp7209SpkLHtW2OcE6owbadBkObD6DF2Kclybc+PQiAUdgkhl
Fq18wATSS1+K5PpcFpuRbr8hlZwdN2LLN+9YaRcL7W03QfcvRuYe4zS5zg1atfXC/UAo1oyq5Qo5
glqZExcdHyYrUu3BD+QgH5x6WYbLi0bKs+tASAgl8ZBt+U7e0EKt8X9Z96J9XVFSJ4lw/cFiOYnV
YJWB1LxXrQdVCaHOSp1qjX1ueEdJtrKvr7yWfBf3p8EfNiTz1D4C6HuGSzDHOPDiOCPM3hWaN6P5
e0Aw/VQ46ba04W1V3LXi2h20y0x90iHyKDMnLWaHk7Q5fblbM6i0v7SOlyofUSLAIJ7rmlHqEQRv
dPQk9HQIt4MbP8/NmY077KQTPUeEklTM4wUnBMjaydioTwbfI8mll7LVXcbfNeQ4euY6V3sLHXFI
NXhhZgSjkWXlyfBTnD06Bjeri9N0Oa7Ov9WluFdWnWuFAKvH1JiLH3R+haQfQ4UoG5l1LmoXMOMR
jcSUPI10y3tAB+xlCSQ0EhTsiw258r5m6RKIAOSqrYkVvwrhA5w7HIUO4HEYumQ55JIipqNnk+33
oZTrGJSe5I/0lUTtApzuzc/ytrB/hNLlIYO0+Vl5sHtKtK7BZp2KWmJVwGUnAWVzATeYKJ+D3SuY
CirgN3NWNtuh0pZoWYX6uxImIQ1BeRhjgulLfhr1b0gz4Xrf0G1e0Grjmy0OU3iMqanpf5ifo2QL
2SzGKvO/7O12Hs/xi5KaE3P2PAN3MN3GJxfmjF6vZ8GxfAgSiVmBLlUnjiAmrMPpfwoYGkj/zG5G
VMKrMRmBNXyNsMoYGoq0AbibnJp+atuoX/H46rKL8bm6B21pgGzJCpIzAbK5Oq1dtQAoUJQo+9gu
RJUjEGEkNXqWcVRXx4etX4i7Mu5HSNuAfWjBhPXzjfT3eKJ/kESjuXAcDsbBIXW3W+k5gNVer1SF
hmgf37BXMYM0/7GqOQk23K3SdaYoMr3B3opCrTwbO4E8WIsJrbEv/y4J65nNhxfCqMeXM27JIdEG
GxDyFXxKl50Br09NppRoC7HZL/4lpJXCnpGO/L4fqV5Sym62cttqHfrh57gvxgRGzee8q1Ienoh6
mv4VDs/+UPy6gb2kzL+GFFM+3zgxYK3KjJO0GJNC2AxCTaUgJVOL4/5ZUAeTHZkmxccwHA3qgSKd
W3ZHs0MZ8O6r36/rXD5VNmK6SlEvMJxRKa16lEy74p8t2+AavVWOf3WS7DBKLM9Pi9cG9Pitd5jc
L8y6qgQDNmQzoff64h9aHokLSUHeMBjxF9wNq5VO4dSw44bpahsrPRtw7iNXdIP5AlvT5pch8I6K
rR+68P/unV/XzquyonsGZl8wWvYADvLDO5pZcfc0aP6AyUj9dsqu8UB5srb2kXDkQ6sbE5NZaaxG
uRAFLnAB9QuR79HYQliiS65VBDwpOHVCe+HoWHQI4U2HUOxy6Z77TAt9Ls9KFmCr4ZdOjkSKMCdj
jnor/kvbN5hqNJRTE3wWEn3vvpvos04hgYhycYJJSz6wz/IujBb6VBF4Qd4ST62hO9s5RzfSajbJ
N/sUrLUqWPQRKxcOHkv9aC8dWiFWfSwRZyLRDhanTCu2GD0mJWu0lHuRQ6Hs2hOE6qBemz5DEKw0
d6c34RolZTp0fEqQ50qionIqTKIviddDZEtjXpI5POPvcvrVFHQ0ol9wG01u9Zcmkd8st1gSoHOf
PPR48xf3DNpPIgkg3xbnlk8VDQbBHc0gGl2sqka+yBifiv3XGxEpXs9FAs7Z6GeuWuAiA0fXVNkK
q3iUNcqCTJKqpl6EkdKn/Yvjc5gTLDf8eYYUpscW7MLlFM+UOeXVcufv2sb38W9NOrJZFm0cd7+M
uI4eHm7Ie+CtfaAa2OV03TN6WMW63ZLy3Yilxh2xx+ZLi+dWQd93LUMBcu2ZK0UlTI7eBT+mpNoO
a2kswEz/D9TJoC93ajhojbxdVUMe3oBXZvfFdDlqUKa0rQwlFYQXbG9I4Sqr1QPigSb55LMkGtmV
dJvhG9328DyIiQtrtiD3grt3o0rnUmA/qfCL9mC9nQc8Tn3JqtZx8lDanqLZyP2VKYlEnCT/m3wq
GoRdStnRPPz4/IQhJvC01KxRZtRf97sEh3GnNp31Fr/hSwohwDZwiiX4kFnx/N1CDTwnym9nlizP
e4tPQ/0dAWIrT16riJU/GOVghpDx15ImHLjUA9t60SOz1ryYcxZCYndIvP2pL52nr8xfmFQpOkTe
j2P2VatiC0w5Nw1ix2bSxVtBskM67zLS0GyTAkCenk+zAIfRzAFDdAF2tPmFCrkvztn/+Fl5tNbW
5XnLi30m2/yTrLuRk6BKjtveKrYQVto2cHpUZex5o3Z79YiUNKJQ8+emoFlep2ys8BZwznOtirTZ
3+CpoY22PdqNH8+Bk2h/nNhKOrYrzwuCbzWUCy++jX4QgFjO2H/plPcgbLMeDi2laQpbUH330uD3
B/QagIZcSYsuai0F1BmOhCzwktQGMddfMTdzo+3ZYK553h8qiT/2KHURzTUomBw8UKJu47FymPGt
JirSKu5njvQ6k/Bc3UrDh9N9i5iKTzJrOrVTWd7Whd1x5opb8sxYnJI2U+PImB5dejtf3f5DNHMw
dO+hGHFEFxddXDg915E0lY5jcnT5jttVUeHiMzsaZJlhHnGmZoT0njMzt4FVox9uEWi8MXGkxJpb
Lv0eRCAHsylAzIWa5bQiADo+irfFvpDJuzHVAvcNXPvE3MiWeyF0tznSuET0ZvpZFgh97VldQzzi
Bq8B1WxUJDirj3HaLhNVSStg/Q+vp8QIMPyqbKRxmX74YQ456sSYVxIYNX/klS/NySYchEov/Ul5
h8MPg2Ll5ecfToUaOTh5FWYvT2KVcQidokTBsJDOscwmiKyf74jp0+DVDgcUNxmXwzMb/096NPjC
a2yMMiIUSqVnHqF4lcamzIc8RNutP9FsPyP8vmqyyhUWTo0DYYC3C1BtISYAXTUNLCQvMm3cvJmp
3Bg4bzCM30GSvNXKEVKst2LryugtmfN9QWp7d/DyjNYmgGk4ZF/g3gRES0lU4w7GyQ45+lyNXZTr
nOTGxXTfSnWGou4ckbNROPtU0waGwIl9rZ5gARkFb1FbrPDWOHcfcBCKcYRDkDJWPe1FdfQ8LP3D
mGGQy9bUCaIB2olypgroBYHdb9WMxadNZP3FOhIS0Qe6ymSbqMxUSLwnjiHO0jvJcqSwppXV06VR
VUj91RRJagGo+97KgnWfKWkv4dFdIaUwUZnVfcIt7+PO5LYU+QsuSUJkIjTGR09jKycYB1OOo4I1
/00J3qEO5xbSdN8E5T32JYQ7KygxTa5yUQgGVHUjPsVTuyQjyLfJk2Oj4LsdkGLNuoPGsKTuLUl9
A2anpAoB2y0Ttk2hjknzLDn/Wcj2TdS3XFqWS/BZhFdF8kvj7FXtp5fU0jT87gHkKI7aRShGuXqa
sM4HcBF5lPrDvY9yDLmYnxqUopAHT754JCI6gkrETuf4Q8scQ4ylkTvENc2JNl2pvxBOGykQvPyZ
HJ9DloCG1FFLmmomKGbOJiWrnhdbPf30wV6/+FohtAuOuxsgPMRXmtLyYr7dyDNykiqvea1HlKux
404IzLS0gZK7eJ+bs/lYfWQILMYrEctOrLLWYYsVAKA+PYeHtPy0yQ7PaASDRsw9PQauGWaWmCRb
WjAXRPyyenbfvUJhcnDkYn9PmFu0x6jRLzQebE40xy/BDWhnJZKjjhloaQ1GWWicSND60zZuBGYo
mMT4PRGGO4WEfFiQ6pitBGE4x5v/vcHoAi31oR6X0Mr43GSdEUChOy/7BdZ2p0N9z9DmVEtsdUGT
jv0YAYs4DteP89P7LewmSaj3iHdfQp1xUsbhzBwfA0Z0rschPBSkXd9k+SiWt/PJ+pgbYbHRUeWq
m1nq0F4+uJIzuGqmbfgD8TLRXcAFYac87uI/FnWAPeDAbqXfj7bCiLAJvAazOfzMENJnyk0E6w5E
flAsXJNcGgEMeyFhZ5zn3eXUdaPFvPpiaKNFXrQ356UXSoJeADq1oxwlfSyARCrN3THLfVWDIw6n
VN/j6Dpa3YaJ11XUyhqmVGuTR2haXymznxsP6YEReS71kZl3d2i44FoIb+qSzqvPMB8E3q3C+/20
n1Rdbbav2wKbEpSiK8VWWBZL04QSXmJIV0pIG8PvVzAMM2jUMr7FIJhek/aMaybyekP5wySEnISS
hzTun2ET3Uceq9Oi0/C0tWUcXYQpRbk+HGajfg1UltsD28DbnzqrQsCi0uv0R2cthSeRbiXrz5ju
Qjg3Feyetec0o/SM5XAsvEyqZDIx9Cq8cBWr9FDMYjLc9mlRkfJMSCyIf19if71hm1A31l2Mjxon
0u4kfppam00RAtmg0Tt4ebFUFbH5RUij9vokUZIFtZcO1dIUeaABPcCXv1Om+TysNrF0O0QEiDVM
iOHz08qXdk3f/U46lXP3pLTpEhtdyBhwFQBaPNw+vJ3ZtOcoRpgublX53isbrUqNhceTF8Rnnlze
lW/Ajgzwd6B5DglMOaNI9GCbPZFfZ+yz7xSKtUctsjPqWSCdzZQVekpPGeUVZXPnwtmEqB9/OUod
OzAjslDBc/r/8xIrHyXnKE4heMY6YfVt1f0IOwOGSjBGBGNQhQDeEMGqISiUxuJSbYoxisBDhRCf
0FkqLJ5w3DfKbTfkAmnCmVN/n++a4J6lV8yHR+P4aGEhQxti+GHOFOnd331m2MlMIjgKmTfvEw7T
narXZ5Yms2jGCgsiZ8WvOqUUHa4swgcTyxVWQLKe+DDPTxd6KOTf5yyrphohDTBFgLB9GFA0pQjO
tvruinOVI8nD5BFI0eA0OxsDwxQIcbIFslc3flvmr+Eaw+WiMtVrq5wB62QVAkV4vdnfKPN9tACt
0LV7znNDBzFjDgNBIbof6Nip8dgOA3mkLh2K1OxWEKFfq1GbqY49rw67hq01gZ/S/duhAFsbxe3/
fcveBw5RVBzRiLgLVJSSuiTB09eGrvoc0i1dRIwVoobHAjQNJsmPRQ7oASxMIw9Y/ieWdrifVgkK
vRAWPuThRjkzHarZo5ZdZdqqbt6G6B8ur3JwEAOd3ossoIzcjwl+h4DdYxo5I6n83u2/JZXsBHgZ
gQWvZWPNP9LkDzA3/07LehrvX0DTu2/yB8o9ZGSTWJOjNqEj3gW7JWS3lTk4I1jCJ4SD1KBkKTLb
MFkYX0wPDyOD2zi7XKDWa4UHZeCu7D2Dg8zO9jqyRsI11wyyiTu1x+eiOT5QKrJZq+Q6RnRJFNxh
e+30m22zpi8MiPVY9/UVCZnaoKOzTG6brb7a/udkp+dMBVam3iQCx6JUarGSjeGZo8fcQhbFxSxr
Ev12jCm90eN0rvwDCKL2nw66sI+zOBvQNFgiri6DeAxpYnGf9HOm6PKyScsxVO31Y7byjJUt6LN+
bJBDCjBu4Nbm58+fv/bpIjThTAq/4+R0NfrJ86I2vN3n0XvXV2Rw2oSlY6auRmehWkeI9cVXPvaT
8FGuhSx135sV71pvTJiQl7Ijc3bIGsLqJhLJyvVcOmBbs3HXYYH9CDLL77EHKJnsKL441i/s9DgW
toeJx4u8QgMku+UUu/e6cqmY0yMBciu7ZVvAxI5VZGUmBl/dgjd+YyfB3xs2sJkEXE2B3b+2SA2U
vamN215uS9QUR9s9E3ufD+qXSAy10pnNwXfizpPeat57WF4MsJzz2dbzC3ljIFCM4MOMHi8aaJYd
/1Q0B9FkKq0qEB/4+N1KLn8GT+nm1FXsJNMwx4VGr7uAsxXx97eMjgenO/ojbF7Y88MyYE5QfyrX
TkYw91Y78IMYY7edwEXqVGG7LqW2CHg8zkLNHMElgTOHSq7y1fvQXeLQYFLiXnlnuERQPFMli+y6
X+khkX8sI62NHAVWgXzO29kREzzoG4iwJNO9/spehMntJCG023B7OTPtdOR0SDhI5urcHBOR1sFb
5zu/sd76qV2lh+G9vswcguIZXHgn+tGtceiHaccQQLEsUlCPSq2HxzqLA9qgdWS56Kg/1eU3DZJf
l2s9GC8krUSsRQbHeXVzYeso4uNb7IQsWi2Rf/99fv7VNqCeju8NtL9z8J6fh7X0ImIDUOcPgqvR
Gln0TWbWAkntJAJWdMKB1JTEETVGRocTOlxeR3ajCcizSeBSKgMgPhPWG7sjFNiN+JnRv1gmz/QV
DgEdf2XMVDIL7Z8mAsiEmCq9nvMAztkYJqlISZtUahe9JMmMdk6b0pbyWYM7cK6sDRcd7Om3Apx0
yaIFWTV4NfVoeJ8agb1WT8K2PZf6pAqF9oIktvkLiVQ/cVtBxlnVa8PfWQDpwWmjImkK7J4pqFtc
tJrZX7+bBVYpfO2ZnNqSEufph9GMHg7I2eQQYCb64r3Jk5Sx03YWIklpsjYWurrCzW33v/pVaOgW
36s/WIXoTD0A/SuT1GgVT+5mFi8Rc4DPRKh7RDmJABMd29sihQ11Cu9PvWdAkU+6n1W9XlRTf9c+
9OS4wRkaQeVpm+38+6uA88RqYFJkQ0KJLcQKWXN/VtnGe76+pO0xA2S6ChsOVap+AffEbkKIg9P4
1V2COEwnDL3NdqJt9r35gDo1x0DRcBJd2JJgdsMYl92GpgUE5LjEd7tgXUY49uq5fYhKYZd9Lr8d
DVaPOHDj71sNQlg+oEB1PrXKOOeRZSsOqscuXG+pRB8AcIjhlejYZXAZXT2iG8JtZNbiJqnwnYQP
DuoIMe0FJBjrt3LHkD4xoG9NIPuzmO7eqVeeaE20f5HKLGTiviXKX4x7qRAo9RP6RGulMw/byGPi
xVk2T5VFj28enK0Agbb0q66IDsxtudUKYv61hZFObDMRIfAjWnEUtXlK2GjVj/BpE7c73Ooct3ei
BjRP9LUo06J/RL2dA2GQwYMFl08vH/JHPcFIouWyYa+SUByBzS6VLjy6Ja1I2Sx45WjUXON/J6AU
ALV1Z20aSThaBTKoKyNiSUJ8W65AHAwFBqOXwxuGOgdV9ufneWGAjnhidQyHEa/xA9skPI72PU/J
/7zxsRc2nOKiWKkgVMig9vNORHFoPwrhWLu5q4YIjeX0/m1eQvkHXO9Q3sk0wMd4E0P5gnD5g05+
jZF5iabUN69nlkKDmKgZKLPYsWo8ANtWvcqMlp/wBm8UBjG0DKI7bHeT8c1CZauRH8zXoJWoB9gX
kn/b/QKKfbaZsd/WSW7bBZ3mmofgS37+qnJ0VJA89gxbrZGK2E/uG8KqVSMN0CEF2KGZru9aSnus
E7RlOwNcpm91RX5K6tTnR9XxRtFLs7dsOFkV+ae65e7gEmytabaZKZ1jAD5O+Gszgrjt3HcKVzIr
8j0avqafKXWp/fdkUPjXAXn6aP+dszzvtXQ5pieGLtUSV6ccb/bofDvINx1PM0arkRigyU3O/oZP
T659apxVmFLTpzoGVxs864j+Qi1SNgnmNADHIDcg7eypbMQzyo97mEUPTjk82qyIZ9Z4jmDIpFfh
yGjZkgIi//iknP+iiphNIDhpgQCmoWuuQkNzOz0syiOKoAkp7tJn0e52dX35bx2q8VMgiRXlI/EN
6OIVXlI+EpGVtDwcgo2wNttkf8Nk9jWgDslnqOGP1XUDGZbgTeLFcqugSAq9/W4zBgBAf63PiMq3
vYxbbT2ovqT4rWR11fd3E28DE7rqXYFIuXRGi+AYOt7qJlDmitrGhDn12FpJVim8xVuBsxlhnPUQ
fVF4Z4Cdph6pQIbxHXb8u+tCfE9YuS1ngeTo7SaW1lGV0mkITOxyudXw4CAxiW0OBX5mwXVRsGf+
D53H4c2J+wLG/Wjy/gy8Dif0YJYB4NDDogWzsSnkTZK/9KPaI8ILMAuUYkpAJIwSIajchtG7IXB1
pKvFdCZwjMm+4PR2hvvhOKZ6m7ZV38jGq7KoCeqedSSVQE1xhIFfA2u2YAkb6rgia4F6TAWcQ6RM
x35FgrVsqKq6bqW8MSaqWYkii5CGpDvw2tUrZB0acnysn7ubKXkLnSNMMkOvrXi9BbvbS01JSMvT
viyWmGgRRMkVhBdJKaVow1syD8PpEOQjX9EMZ9nnssT1IZCM1Yk4dm6feNLFSl+hULe0wdEDD95s
Zv3Zf/rQHmgnh3klGTOIEVdtRH/KBgg5SyWrdfa5Xnmys7sFtq+HQ5kaz6TbD+Ig4OKE+AD2iTLh
uLiGUXe2vwsbizO/neh3tgtXSJniebl5A5XaacMeEl2d9wl9ruRzifdojNirFH4vVA2Td/5Omk/F
xA/s7EjYAPSOwPRYF5bDKdCuhKle4jcmaVDJaFK7k6bqRJ0DdPPEZCKu0SPGVuMPaAO5WkzASUqJ
rG+OpTVuaqka7/qiWuglWs+KxjI70hjRJCkb6PGgbwGc+lS8Lh7W7/+K1hozqjfZxnXLh4lV8HSC
h86E3evbegLf1JJ4YgcarTzDJFTx2NS+Z9RL8k3O4aL6kKuHYyiKajpG7SrpneeeR2qktAQ+t3zK
rPFkuao+pzPBJ0q5safJZCCuFBsFR7BclhuR8oE+vGJ89UK4Ja6dfsowQCCRIkCH4ptZKA2P1ors
8fVjm30LAYA4Q21AcF2OcXiToCowEPqkJXvrvs8CKSP60hYkIYEsEHH90fMj2MXNzXjAV9mWxs+l
txoriofT4MCzTz7uDmQ3O8odyoFgefLRACeYMPyuHAE1urV8uzgC/eXzbAwGzCsvS3a7hlJgJ3Pq
rXzURoMCBD0D6yK60HfMQqqAxkho36FZRiz0zA40mVf+5MvT8p1xfixSs7gdD/2t2Av3Mp8CF8na
7T//RGStb7j6Tx+1KDD/2O1cJijvGhM5hz4Vm4wDLxB4COT9cFg6PxBiVoRjmywzxbJKJ65zB3Ct
PNs8jv2+yb2gpQJUISD9HAE3JJ3ZyK2Fs3gOqHzJosPu882Ei0lb079eTOx55QeAzPDLYicqUTLM
2K5nOrJ5YYB5JYTw0wXBhh7K8FiSk+ffh3auyzZ+zqitZ2eAZWPFREyFC7aThVQMHNTFsnO7gDQK
VVjLeW/JnHb8wONLI0/hnSNKtgQyQbWY3UFYhgsuPl+3fVfoNXQpgprRm6bLz2pv4TSZN5jh8yIa
cyuG/AtSi/TIOJsYqeUn7sAYeS3SJbWkN8px9+3Dd90o5KtCsjHusgxIY89rByX29OYEZK+lJ4gI
LVqeMzF+YhOpwPiuxpAzgWQAVDrwaaSwoN03wYTihi1G8FVRjdaOIw5O5ei2PxtZ7JBWhP2x9Mhi
DOcs1kkirhcPxVeJLw/2o1Abz+mJS2+s0AB0I5+N7HoH+YlhLutsKUp+HNtZtJ/Iyyys4gOiTZBg
p8u0IgN8b9UYSs1+99HimhPY+F8Abe9IVdY0bKUmfEcPFt5YMtpFr7p5XNpkewBs0517p1FBywCt
ETmce41inZwyoOMZozZw+13rx4MIqmmpR627ILZAhjV8e7Cljf3mQn4SLSCpvoZf6u1KjQueL9fa
F5WM3ulC121WQ4Wfz6+HrpY4WLDAdnBhoEJf+HskJ471uq+5rhmRo6YGjWBnzWjDBg+LKwWnn83r
+oQQStY9gV4ITbuufDW7yGSUZVlBw7+lReFR+pFGCUiqEBe1xcOHLcmLWDva8vUbSXPtOXFi9xYN
wzPVDK598Okpq6O8KMyyL3HCa1kecFIKS0PlmVIvj+coSI95tzvS9Tc9pJkFzQF0fJuiK5WNar7L
MO5c+2myTHnZH5Iq7m6q8IVQC7KypFgGtsv0CEsGAPb7uiwenJEgSDQ3vF8uV3mzU5b6ZIN8r6bN
hotBBiYkQjnYW+avLdkG6ludFqNE9VGNaYLRGEiU1yYRk0pjf/coQjP0CoMlifnYwmDQ9sR1hycJ
ZYbb+cWzFJYARh5UkAobjMivSjpVfmWV4rd9gURQelWZbNOVQKTIliTR8X1VH5Wmu36d/8pu63xP
rOtqN5pQUUqwYv2x1dmho4POZArh6tpOKzQx/R+kH79Vde2CF4a7SHTE1VHiWVerAJeZPKmIKQOa
nYw+4nD/zB5I1KtNTQ2DFmQ0rAVHJV437qsQG0dCWINOhVWc424cTwX+e7q824aEZD5Jp+YfiDj1
HnqhawD0wj76G/OiQ8Ogz07ECyZdWOfH8T1qfDV43dcjD/stGu16J80FmaIY3ttjEb9jc9lcEUXM
0YjC2nSe3J6BtvNJ6KSDOXBaxf61q8clPXrqzJsTsdVqPld7a4Pu+/Nf+kHiSxMW6gOptxJPZC4z
Vy0IKbhwjRi2obGeXm8GnZcgnD7ml1JpzKzZ2sXlHAWQIuHx0c4URJAMB9g5/bFff/MSn9WCkxmo
82MYXeS03iZxGIMhPa54D8NwWd1jDhUFuONZ6//L73MDx03CmlRV9twSFn1e6j8fRLQl6GL8QNMN
RoRCQ7Ef25nfz3gvpzcokY4fKbrXxTsPE7TfDD0FGazimAXiUlKct9V00z0QcyNH1tavpNIwxPYe
8SyYi9W88P6GbwS8cNy34zBYi9ZfzVFtMS8WVOitNwH0MbTX8NRObLgtu2Nxr+x/Xr+WOxVwvwZ+
9lB2WD3QvlelGTpmj54rPBEzI2fdGvlGR6YR9nDdkfpDDVW3pwrUdkdYOkzWVvWzUj+tUb30BSgI
GSBWlu4Qe3x+1q11blwCQh/r+X0wj1lWckzmHYDmZ7KQ6WA2iCAMwC98iX8Zim+GROEq2CgqQSg5
B0QkE77+SwBOh4MGZqcYujSUkt/2cjVYsEOaHJGivQ8E1WihdSgOls6QW0d6jQByiSVH+BPvRotO
sLfCUHKH4PxDqTKzaCnAQY7cYdPBzoFH5pYuTXvF0IJ1yxA1ZffkLP0QxPIGu142R/LTG3W0O/Zv
z7BsNsEKldlgcB97SE72og5iaYIvqVDzv6Y5Fz12q6eSDSzKOQT0FkfY+iP1GRSZ7ifUKLpKVzMV
dCarTkOQ9MpX1dZj2TgCrg/GMwkpx9jo2eN3sAKK0SqYP30EmeGrHzDn4ohUeS8YgvfiYXB4gDGe
xMqeHKuQXVr5Ea6+kq5ZvrS8MKNW8K5JW4R/bV2chx6yaIvQBTuDrWdUE2lSMcZjektfyMawDulb
RxEe6UjOrPvCkWgR6g6RbMTWGDcIZlSexC9DNT7YCj9n4hwW4t2gza4eTYqbpypl3UsewHvXaHEM
z68AivBzXCeUz/9hkC7qniiSIoZisAiDWWwKwJIULnIaYnYz1Cf1IemPL8vsO19F3WSXRmNwJD3p
yN3D1OywOXuIx2Ab50HlHmndJOmZPbsxtcdMOcAv71FHxtdi2y7aMqmV56noaNnuU1SHUyTzXpYM
6zpI3Ziy0dJNtycTPsJu+M68o029hbQQNK3Lc9wugUH03cVd/73h1K8yJvUq0vhZSI5jyHKV3i5D
/SF2/bDh7r38CG2sjzfrjtEKI9tq2RWyptuclE0mk25oJQFQI7LAKtWEdu1G9mFlEj5p8N98flXZ
1mxVi9Xu6cv6G4fPNkG3YZNCDISh0F39TNn8/Jm8IgdTfXImDTRuWVEeUMkeG8y8DaIZfF/QRhlO
LniZlJsCk5GJ3T9olJ8bUpjSMzSndl4xuJjbZegPOO+kJQ1ckNF+OtWW0EGcyDSiO3fpy0d4gAXN
mYU2dfCN3ntucLkbpF2hw9GO3w17K+ekS+Oq4X0l0I6me5QgAp0YtjYmoDfH0dEmTSNzSBWqXmCG
7Eyq1idedg12Fiy0oJ32LNMnoWG9Otf4KYnxQjlxTCOSwPF3RQNA50bkAxU9Jm0jghuIdXrFLCy8
1F/LU6BOYmzBkYRZMHzbJZqaKyspki6TjUTmKe+nCSqje2kNQnjcqtEj5bK7FsdiNjDZcCO2Y9cY
f4lNM8qz8U6wo6Zz80LGqtsOQOGgYtuwloeUMKHhi0a1VWFczZeRIfdjNfhjNwPjXDUzWj2rurA2
+VBWoKBEm9HMqdOIRkLmPJhMW9QoEtv3g+4LqKb/nZ4hGzBl1/EZjdIyl0PpDRul5A9Y+fKtSA8H
In6CamsUHXGh5dlkvqWtcqot/PAT7trMZSTc+Equ+jP+uWm2BG8PO4bfXpkE6IqHUwRqK8DEyFZJ
wKXUQxYW1+5XPtmxiBcGeazxAccLf38oylfLf3oQoOcu+hRzSPVNEO9G/I9xH4bJ6J2WsTjlKJYV
F7Jbx5H1Ya2x7plVWTadweeSoW1snghIjzmgzmlUlPWon+/irghVn4nP00U0Q/mXRs1UUUpjCQg2
gsMZwhAqjLm1fxGGeYEI+ZZ5ElrdmokFq9izqp4xPTvh1ka0vo3rldZwP4UnwHn3WtngWB4PPkZp
PlKm3dXFB++jpxzAiuu1iTOLgqwtGU2LamH+F1OIr2JO+0qzfWYOQAYAB4/1espjZnHqn8fEAEzo
FWokZEbMhojRUE49aJFn5SlmoFTergLHl0giYIRlkwtNyOqO0IPL89+sw9Rh6jjW8T0dRHkaTyfB
vrrhWH7YImeHKaFXXiarjinmsnOMl1TipFaUB8Y0ttw2l8H9rLOKsprkd72F0TgBoJKLFgSpqwgk
9gfK4m/FvNqaBf6NGIp2rNkEC0FxV0FQiwYIKLqXeFK0r+VW+nL5jsHEq/N2h5Vc2wT+Br3I665d
af13EUWazEHG6CLLTzxlCe0+QRKR6HtohusBggo288a4ydCrdv4toHHvL4o3xjoTksTOwpjtbn+p
i1ZnIMSIWf5UHV3BcIxTtYB8+T77k+U9inpIO0ftBj4vcJbHD5XJ76OVSKAxSjboM0ZEpfrII4ST
QmW2MwXRTjRQSxj4Fbi3AxtFAEgCA7eIaYh1tlsSwEompwybKZqDBKZzxSMZ4kOohXmDJR2ury33
n1b305YLczqa+JOQ+DKQETahjSpnMI8UYQASPjjzxCcpvSSG2eo9WLYigruFgE+UyBovls0I1YyR
EVQYFGDZjcJIHsdfIPyttxIL5MlRN7/Zk4Mdk3Us89CMHfKiU9RUOSFRqoN++E2Xs/pCttzfetnK
4MTf6LrksWmfI0/8giNFd7ubTR8uGUZBixG6twtPyRYyLx5HcO7xSkUmRn2+SfV9xat+bEYB3B0w
3UfJmsmvmENXoDIhUqitPPD6C2hgP2mFpTGpfoJpTvIbAPzCYtDrLWEfHMgZOj9KSuTss643Iu5Y
wIK58Q+TEfUVxrBoEN+v0FuHAwq1aPcG4V3KZGnG0WGhZm7zxmNVBd72DIOEFk+/CGJSMpa00xd/
x9p3uJPcswHiOB/q9oKFJUli4tcP+wVTPIRz+gSXpnkKDy5XsD1D36JT8oKGNsuirt/QHrExzwLo
1ecP+Y35AXgeIOT7J/mSJMr5WbktUKW7cAioZ8uctJz8WAi9+DNJ6fllrruzEMJ0dTX0UMWxUKDL
vfXFWvHAhviVInxuJ353th2B187uSsH76fi7lF5+TVdUfmaedPYoukDwKFAbp66J2RfwNBLkZBaH
rqUhaXj8VayLm6wK7DPGTARkr4sF39OMzApA26G8UK7x1n7YJrbHYyiAgt/blwICYa952f1Rpdnx
YfBOTKbRQ86zLD6AwHupX0vO1GG1jirqEpdEjUk99Z5V8HYdusn3eV6KCOvpXWLa4nksXr/EoQ0h
waHZ0TUMihNz3tqQ2JEGxQwgn3nigJu+b1zkmq0ZxURpvqSawq0pvQ+ZPLRuxzNaVNMtYFn4is8N
/D2CMIPE/UU3Ga2XTCNEnOIH/zKY1PnNqQvLHwstyYqpbaoy+wrlZ89rlh+eWa89fg2lJojENUj4
gc3tR8Seq+1rP8ejULNYejBm9rRENr72yH6HJ3oUR0VmErAtxU/QpdqGm0ZcC/mt6XTQfD3XiLWV
ua1Sp7ofbtT9gBlZwT06Cpr1Osz81zAPH4lyPJfsBZvk4Lf2ZdRJegcyKYPgsiX89QRxx+2+YHPq
lc6Cr519uz1LT4jvtvP+VuYmItjchwvfC9qhjlRxK0/oGct6eOW57gxDsa0kGW0jGr1Ri196pQTv
oxCEDUcGT8a9AUneqzDEzj4UgUjVOQpX5UtZ3lDaq05VRFKZfWP9bbn42VbJxJe8G3sEFHZ16+76
1yL7QyPZjal4FhYjhY+Qe4H/W5YYlvCPY99DMyAJdIJ0mIyDwpzAaTeE7JbnaAeRui05lFwsaJOK
1wUxXf6Ce+9oJqo3k2Z4a1gatYJk3NNjAu1iBx0HTB4tdThmuxyGncF1+wix5B51uK7eNVGnVro1
baIIGQ1JfrYFUJskj1amJcDwzi/oeBtS7FsFtEg8HPkyBJL4VdFcaS8G7ReYlZFkfgIjjzjyjf9O
fjkjO4TivTucEf4e0esGhlHqB01B/dD2L1RT9PO1gddz0XEPRS3Na2fPK1sKtn/Ldofm/iOVYMnA
j5oc9PGMPwk24TrpYwXnE3AFU1gg+lLUm/gIIm6RQqtNvML2Rl7rQxI6dQ4ra1P/1jzY+sRUrQYq
qX7UYSdzPlvVFwgs/ytLegSqAy6QSAC3q8ifHYWutadnmlfi3l//upJcL9W+oXLH2jQA9T7BK6H/
E+UX6qHEUCQXWP03Cm8UZoTcmej9lOqQZxwiDNPol2DLeAyIE/C5EEJ8bXiUzEcf8nOoStVj2fu7
9+2053Lwg1DLde6KQfIUaj6r6CHkwLjdMofyTT0kEOunYP1bl9Jsjnr03nfxhwVZEfRv6v1IfbCF
2zDmxTMqrhmEmmuX7zH/i4ugkfCPY+5W2JZZIm+6QbHMbQK1ZnrKM2jd+lKkpAVSo7vA/aJB/be+
slNwqHdoi1TJzipyLfBtW794DVyAvPSNtYqs2U8KE+o9dKl2Ai0EBte3WT4E9j+WJ8VcrmWSfHuE
E6OzIXs90+0Fg9lw4msxBdpmTOmuwqxUvh6mc136YP0tRuum1kurOxAqPmkx8Dvk2p0RqOlqPb1H
ky+p8IF4vKgVCT85EqItC8nRVbpt5S5f2S0PxZVRuX+pkaKG03sg/f12JR77PJ1xlXMEoTKTdQ48
yyuyE035KoiEnme63zkdsfQsx+ffWrVTmsdc+EA1qhaFeN8oAOhcuIC1IWhr1trbuoau8lhb6hN6
rX1T9VBUGhbgmqPmIdB5blUlVNQLTMA3AzNYstsFXVscCd/9banMGAMJYyxhbkGxd1W5MjntagZb
PtMSlQ3OjpgnSnVQ9N8nJoI1r8cV++wsEFHQaTCsQTzpzeF1HrHpgW6V5Pg3DGA0Sv6jDUQnilFG
qZe/aOFUQ3VQxHFuVOvvXSPLfh3E/z24exsTTUKaRrzN01rDWaSObhi8FbjUTRLS3fomA3JaLk/p
ViRefqPawhdwAwIDIRJzdaaziE/QXE+KNYTg1cfqZ7xNOOtRlS1NDUbKZelwYMAfKr+X5YQeTTIp
cvei4qlvLiz/qToVKCANEic4GfzEozJz9Pica514wEL/ay4vnbjrbNp6B0Z93uYb1pFwMagIkg+s
iE1HWWQYuIkow1uUa61I/MV+y/R+e7PIu1VaYRVdQ1GAq++yOhJ3zxLwKByno8WEbXNH9SdWdhg9
IDxOouZMAf74zHaiIFe7MPnvuDCtm1D+WGY70hsKo0oLMKtz64+1hMLPr4YyXfk9K1fxHd5beICC
vd8Qjx21AOBfZystrGhn8j0EccQIogX9XMY0DM/SdLcoN7qMbp1uZop25Iw59lr4chYZSVsESA4G
7wKiVsY+R5tycmlZDKie8vcyH+SweOrrX4FrRsKlVCS9v21BISdDVXoZ9g+484lzJFKD+jDgjDtH
NtqEVkLI8bfIswtGfxrXiTwaJ/EzoSi2dYlW9qTS0kwkYE5mwTp1Sv4hyKlkspPB8IIT0sOMYEr8
gf1SkleAMRcdSUuTdzWhXM9AWCjCitaglELpdlyOKxQ2mkHbUY9HU4xU8Tm6Y7svSHy+uLyn1FAg
hEjn+h4yq+Zmfs4kII1dKcI/nQfQofnco6lIDyKkt0v/2d/hussdoeEegww+rxKB0DZPSfDKM5O+
RSmzfqlEdEJTtFwQFZuZr0c91d9iACUe0e7Py5q4ZxE+PEGqYj37jiESKPAttmL96NnNvX1O3lRD
fvs7lCUxxcjbBZUy97VIaLfCkUB6JJA330QeLyEBivfWMy0F2bqxJsAy7Ezfy61YVmPibMSby7Bb
RUWd7+FmfHcDHm5+Vq30I8U/FA/giWEX5y/hEaRr1XHadGZd7wBuvLrYEkWomiWfbkDXVvST/w1Y
8xTjCR4jZfPFHlBG0CnyLqQ4eiN7I6Nr88VZ1BId3/woGaWEBJlZQn0BgYkENAEGf7zOClLlFUy0
UMbPOFk+nLKyQRhw2kjxEe6DWXfjLjX6BD9sbyQDuCJxlC0oLEdWtt9fyDfQOZZh72BIjWLTtzhJ
+HDCrTEWZ0uJdJqiXxmkbv0LkBOKZTz5cvSZCqWBZdRFECAArltkDnnDgn3nfjs/37FHHUQNIHza
tODZVE5ca3KB+0hqbZoN5rlgb1whAso/DWu44IJBVAABKWZuY5forTioAjYJNgJ+8OVuHyQukIsJ
jVCgMl5CoWxve0aIhaDnnyLawTG7tkKH8uIMLLhMeVdRuc3LFIJ6vcebXLKy5jg1XagVgClG+Mos
MvqtVw2OtS9Yq0Gz/cownw2r48nsFWwZM70lyPyrmNzdLB9Dk+Z3jJN1AlyCNqM16+aaBFHRKsps
nP/1GEXOtIioM4iwejEU53wPAUCTGzlhjbnhfWLH/FbNlOtHkNl22gSlqzIFNgOh5VnVbwm701En
kyz61NAJTgdrBTBPz+Ybzpdo+9LBisoNOPPuiqW6QJGDIu4AR/uuKiitT4yoHg71NlohS1ocejyX
VHPug2zhGspMwmzUTlQTFimz+L7pX1Sah85kvoWnYaPxkLEMSxSxCdJ9cB1klgELsTEuXZ4Q7a5F
7SunwcJ5JjeiAGFLnpYIKIGubdyOcXBAL9Dcsqg8doJDwqzsQhaVzRt7cb+x7rTudJzXA3wgGHtb
5RjTH4bYGBKoPl1FaqHwhpn2qfzAyGJK/R+SomdE/KJTlPuvIHDODsgyVZGnlE4/dWsQ8glVbaby
+us70FaJLTO6pMrg9Dhx0Q6LKqICqKcFVANlgCKn/vAaLze/b094UG0IgWHmZe9SANJwRQmlJD9P
iaVE5Y2Jw8hsPezrsyH2XqF4Fj/6I/NCjOsBuFH/5eayOBtweOythsscfpWWsAUPc49bxHXDGm52
nyI6JrZdI4OC6u635Bctf6UFrv77j3mgRPw9RlvXh6eEZNcRSDSHqn4SzkYZjb9e5xjjvSxdXgRq
APgzvpClIvM2baTcssWnKzbXVjzLVphPlWwGKMJLOvto1VY+13pLWi1BccbQabdCkaasJTkBh67t
tdFAUk9tUKbnLh68k9SPOPn6HUQNBR1qDj5UIEdoVEbXeBk28WmuUbgMNOfY187Vfuj+ADjXoP1/
KN9yGmu0LyENr7ely7upUsN/bC1j2MbgaDTEJUhpoW6NVa9V3TEIT5W1YwoL+1o0/Ik8MuAZt85t
KmCXD11BHRzrHkCDnI51yqy9Ig7q70yF2exKGGeWbb5414wjmZpDx5X9Sj0ao4C+8ogaRpHmBTa5
5jlJwzSpjcY7zcps8kyM16kP5IeOjIcxF6fWBcIATXYp2QsyVamhOHzd92+sx6IkmDsCXqU+w6+L
OtOTwAtQHU1Xyk8Clmlvf/klHlkTHjNzNLinsGxwoJvOsHbylrUKw+7xQHN+c+y6zFm9lsDIKFiS
7mfQWJ/r4SdPhbpVMbRCtEaRr1hLmbOGvS00IPIbd/hEbQmSBbUQlengsNDFaMDr6DdDvaMWa0hX
KekYHcF/D9TqfJNqp/hI1oYetnud//S70zOAatkimbrJ4Wy8OOf343pGyCJaF7lkkCqaAvZj4Rr2
UX7x1UQhjOFeLoj/GwLdz/RCXpjliKzZvjYsJpw1MBxVY/sbyqgxU1hTcC23wojTwWsLYaG8nvzb
vjOH/xeVHlNC3RnfASLjKdSl9fKIO+nY2ogIs6iJ0/GjnBEAAMdVHpljqeCJvorhS2MZOIEmszho
V/Hf0I1sgQOBAmJeDq9wNFFbfUf/+VT2dFGD0i++emM0AmaCyPwM03D3ndWZPBHrl2zyb5Jb1D/Q
OnNrZmh4nrEW7qaoLND7FvVo6vI3W019jvGHnmAROjZVdK83Mfv5AcXfZ1xm8AeBikJfuwjXnrcx
VRB2dn+1L0qSum+0ltG7vxqap+BZOQFFDofKtbhnMDRb2CLHb0PhQqGMxEUjdxoY4X0XDDhkSxA6
pRUnYrBbGJqw6dZtij9G74/w2ZE3zoFUAiKVZQSx9vg04kY8hXzXojd/GhU4SwUlDG1SP4uTEqZ9
m1LHcP58i5F5jeib2Dx/Goe8X9o4UrHUp/XZoiDi9E+3cWyhbhof78Sctf0p86Pp73AQ3ksGMklO
jgDovk/Zpto5J4enYTeZgMty5d4VdMCF/dyGUlY2v/dLN/WwUsVS3bDmEDhz+sFSzhKUIE9KQesa
8dCAZ6E9wtwm74FfGc349jy9D8ys26GtTMbTKHvXO1wAF96piZaeYjzWhbCEPdDo34U7qY7PuFip
AaLi65bD1Aq5pmejFfg/92rM9kSsWITx70/1Ke6OQcXvxr3JylM+/vkL9FkueZp+R9XRyxkIFy1i
CHirhNAvSx2XoyYMYd2Xj9QXTUE7c2o15lVZ7x42teN/G8QAQfP2dhU0aLR08ryQOCcTDkTU9Bva
A8TylP8DGWXUFSp3mqS9N/x/lRDPBz4/KWdOsTUotNl4vzLPn4mLHXDCOO5T7ZgQRS96qEsUvAgl
DOJADZRheLlpjq/11OnsvLbjQGs9GkRDMBjQkmYqOLLRNwR9RtINmVNf7qLOPIajYOF5BUctq/ZO
9b9c9qsPV+OcjF/QDHPuJF2HhKuuvLGfiEQS0qLP9bZWnil3ghsLlqMMJGxjc/c8dT8anNNOrpYZ
A6OxLi1xhQfV/A73vdWuoj2Sh9XrNAEUcb9g9aJP0lXTgDja/5AZiK8h5UZw2FX/p8FX+MeWmbdI
nrkZgg5fvSJhF2eFZnyveWkVQobk5rVQJtlixYkNLFIH4ldMzgLkpLWlXK6wPlBehblnu3qSHX3w
GowMHr1dKSuHuWKWX6mGDGv3ZI5izJ72c1n6p2zgXUp+/Cv3wYGMRoyoZNNSxR8lliA38nsFnggW
WJGdtm5CJhTLI8r3ikk33QorwqnBwDodCqZ6QHlh9BxYiFukWxnTcuqzjO6KmAHgpWbRan7238p5
FxwDk8YoFZh4EAtG3T89IhzE50mwOGdrkn3heO45Vnyi738C46KSMsTVvfD72CQOYPVG3l+RJmAG
L0/Ev129mouCoNS/7vgujdlIrXTxTTlKQCMkqds0PqHjEJoaKbs1Xedq8qpzhxKixP6QT388Wxp0
aaNeN7nNGpjMfiiffYczPKlJ81uzz7OiXr8WRq5wj4s3SLJeMpP8WEVM5oB8zrvdlubNDiJcI7pD
aSXkuk04GhtFwFLW+YW5CRqdF7sarAcmtLAoSZN8y5UhVHV+c8iLupXoxb+kKsGnH0kcZi0FaFGy
8LJs1zKpiFSeifr2oNDi9hKpc7RWAHGivKJlznrgS2ShHtNzeJIChqkYqBaDIlN32SjMTt41JuCg
cEYODt0OcJ8MS34AbwuMA7EaV813npwnMEaexh3QKXb+EUIxNcE9366vrMqnRfQxJO27XcGn7rIj
zE/gid1VpxApeHRD/TQk6yfVHao6+MgyZLJST4/+eebRqPwkl14Ti9jm5ItoLn+TrapJyH16UHVY
rPIUWLTdtd0APaWK04vVndNk/ItMJt2ANCEWFy4/jV7bgM2id0xIiX0YNcllcdKyV+oX4vfsiVsq
mGjUQDih8gtXy0nspHdRoLqzYL2/YmC22CHOuUsfxwPHqcJcqsbg3xh2QAXc76guOpDHbJ62iCxj
/ON5zH0qFtTlBNZHjR4WctgT8IKJ+ZAFo2O7W8ftYO41haVFQv5Ia6PacSZW7IhJaRz9G4EupTn3
WaS4e7X5uvoxLfYFTVBYyyFPPYZHqV0G4lWDDzYAPN2Iz+/HRLflOFv+/Ts0qBlgr3TY/W+s7xKg
AM3zExz2JSWR5zAeNbjh+XAf6gc4bQgJvQjGVK6J+hFbNgpXuTzx4gTOiHH34XtSeEvImRoN4KCH
2OJDR+svv86PMAW6OZ25bCt6Sg12xQHtL6f2DBjZ3fUdRXRyJEKc69nmU3e1RwKJOwZSaoZkqThR
ozDb/lSJ6FcUcYVqocC2r1u9T+xAxafUCzprwT4LvVZO+jh5mVoRnC98moiZW+PKr2AOWW5AThKw
8lnwPpGstQBrIw6xsOdqGee1wLCfg4pZA/d8PEthtdavrjwKYR06W5M5zPyq8JXSTPmnn7zz2DE2
YGgSKJy19ATk3GHpSpKTtCaWRavAL9UKRUPIpwUUA9IKp78/zP/f4JYrB8YIGd0udseeiRwP+ROz
NWOHQGHtvqe/jOLTHeeMTpyun17lW2iS7Ui5MDQlnTIjLjJ6MOVoagpifkskawhRO3/ok63aHr9h
boqT0Reed/ktaS+FEUPnP4hsMAl4tz8Th4sKVWPS5NXw+V0zEkUU4MUnJZ1SQph0FG+4jvHC2x+l
GpHXsrq+qnI2hUF5YQ1fY9jTMhC/+bLawqWB2fu4VJjNkWc4AJd/FEUCu9IQZASM7ZtHPJOw/e1K
7oXp1x2lWuYDFzIF3tah/tAATIiLL1sx2fWM687uPwFYLqQaPzFCuuLBqHsJJwfoWXju+4p/r5XE
JKqwh1jR3C77+lKKN3pzMiLGThvVBumpApdQOPkXbUo+IsJv/QdekDXW6WAqh9hMmh4RYt3JDw+e
QEPkPqhzV5ZDKoQ8E4/okoZJ47yvW3htEUGYgqkBO23TyJfZiqofhAelBvXIOHYrF1d15OISiGS+
l5g/xFjlJjoJxxZcfZztwlZCmYMiAuQdx+busVNCNLtIP0RvuAjd9aV3m8ZCIbE9Tlw8hg6Gg5Rb
Dg+pkvT+/BlcoTZex60F8aXOLhCT7fhRu+h7g6bntXRb1G0c+IPWzUE/w3B6F5ITj2eNf7gHHIdR
hXgP2y9pLnIVllho283uCvW+jBO3R9j89u4ah0afqHatywJLAF8gmz54dHPl4PUJKT8R3cVLMbqF
L2v/UgtVxDO/VCI1vkDUo8WsjOwnZmlBVHjQpWo600N8LDDGAQz3bfbdL1JuRnY3RqQSKmNUPaZU
oZ7DOfOGn5SBRFhgyu5+RHGxEeoyoVgn71snMpQkPdiuMmY338oTMEqiy/x+/SRWagahX5GyxgJe
zvq3vMA7Ar2iqTF2cNkFCbkazTQ+PE/s40JYGv/tAop6nVlbAvOI4jnJIPvGSeVuKL98tb6kPvWs
M1EGjYdSlZOmXYGg7QGM43mJ5gufkOuLesEEBYYWm/xDEQZYG1EZdU1N1d1K5lCQW/8A9/9D3qhm
6rxXVuHyqJVuqIoMeOCDpbEntlvlcCoK8n1lzkGAuwjQyFjLm8pxFEbERps1oxRq30gHkoxOAakZ
zbWeucPIYi17HPIPOEJiTZviBV7EaouVTxsGyHNSz7vyD94c1Bbu8vWpBQBGW1sYdS9vmKyElcux
GJsJVp7Dwyrk6Z/19U2aggr4xxZB+ASof9fcSYkEguUEzCH58SikBcTXdhWtfqswGNsGfOyKJC4I
AbZbA7f6gsoxeJtHbi0JsXHDpXZTxaM+WxtYCWY6yB5AHnMjZasXBhOLHI98xJNVjIQkXmFEepcf
4atv0ApVJRyC0fXjnZMZfz/o4NdM5xtAcnibt42sdmbOadXPS/G78T649lJ5n1xXWevJfwa5EhP6
NdN7xkzdhWtaTeT1NncOTs+Wi/Jlv+UPxNLfKPrsKFlYUVNDFH4RWxb6O2wyBs2Lx9l5izLy1gxi
J2uVS158maS8MAgh6XLsL5PTTguCxjDsWbIVcxjbLrM2oJUXdFZGdG9MMvdT91R3gnn1Lopce9GZ
Gny7Ov3vF9k6+PF/E+oK0KmVzQH1C1ohx5urZ4Ret3IcoeLSM9HbMAJtpBa4oAI6nNl19pHii3oR
agEHpaCzLsvnAe4UsWgo23G+JoohEZxTl/XmdNbZ7GIJy+dXg43AOqHU2BZ39/mAevvZrj9pYPWu
s5tI81yLB6W8q2A7JFLf5587GaPerlyhoTaAPVPvdAb2QSTR9G4CXb0dCExouF2vLNFtfhMKubgC
zwvj/jQYsYGLHBm5x6CLIubqJx8+dZiiKWuuBfrAYqIcq9GzdSIIjM82rEP8SJhkgH5QDCbI3t8D
ChF5aV9p28ooUk89dbEt4ymBrDqKfr8X2dLyiGss2g5yyZVf/XtqWyn46tlQUCyJrbvlQUbhSRDJ
fJ/z8nDHrUYb401hx0GF0f3S0Q5j6E69ZLRXzBusMT4itk1ZffwXhInsx5HRqZIE0xbiYidFPJ/u
U8mYAjYaC9cZG/9noeWlT9ASeFNeL0xQktDKSwggmVFbD7YMNSlPQcijKLYk3fodsB51llIP59Jy
rPhoLZ+1irZn/7qJZ5mkGNIZJakIxfuodH3+OnZrh2wwsOjfY6oSjgB9IqdJ3VoxMf0LuigLmIHi
oDkaVHOZXDhmXmniCyZPRspBz729gUAkv1YcTcsqyLISblJdCTNRJFp7VBGPvyCf+rBOXmWUsdoI
YcxUfPRlUrQNhZTYXAPJsEQPPN4mfuF4EFPkvgnHUSOofwvF0nUTQ70pZx5ebZALOvhYoZi0Urh6
dBpcnRVSB9JapbhYOonWl4ToURryQnbd2JIFBJZyrZhEpbndeAUhFvOCv5ysnUufox1hOH36BW+d
aMna5jlgREHteM+vHEIYqn5Wnf2JF8/ueiehFQ6o2hmg7FQMTgZ8MC1v6rd4TD9NQ/PyvmOLs+qn
x/5UenIcCZ9KLNaXvEAiGvwI0rAB8ot1q9U93NErSNnqKkxczB9f6AmLNHZB4+FCBfrdoXu2yKlq
Fu5EKfZcGH9CNLPk26BtkBIPZ3GeJdw/DOu4MHc8ISr8nw74j3m49Z7NSYthCFauF8h34rO4fxcD
mpEjErXBIDpXjQ7aAwTl0MAyuRgF8AHSUPtupqIAGzeU+vKgtPCVvm8JoADkaU/5jeTqV0sSPvEK
ukUqUpTxNqlgiYrwK98Q+e/F5jxOwpkSVERXNWpr4tGl/WwFopp/QHui07zBdp6lzZOjERPf2Vt5
T2f0YX12F4gvuwSPVP/kvqIvPj4mXhJYVRjqHl0PcI27uU5FGmIMBMWM0XDjmXOj8Niz0gNFvmNY
WMPInia7YrRxQhm2zX3ftRef8eXRtqpZxdX4NG448arzUVGxa7k0Z1TWfJrLXDw8jZYa2/i1a0aX
xwayNm0LahVRhmUUbP2hQSDBGLzgG/It87JAG6jl/5WIPrwnKOgoic1b1bRjBv35hVjwhDN2dc6h
qhuEyB78i4YX/fcDHy2DzmHUoX5lcohfpNdAaurylCH0cZojzljexW3/gWB6nECBbqxABgPpZoq8
YonQA4AxACTwdzZhfC96C9XA6DygeKO3IyKKNY8O3d//pzJ1T/lYR+6yWRERpDt+vQTleC95Qf5U
7bKzmChMcoe+LVn92zXeXkyNILS2nwmudGTQZKdLtKCGPuJOVbT+oi2REmlrIPeAtynjUnjEe/dl
lfNj74Lo44y/NAAvxZN8fp3LtBrwCmiNVbzHGGYM62DQJvLQwhuMGSL+av6Hkh1fmjoeon1aNFkx
oGwjmHD4Za1Jr69lY6YaWHL5iRuK3rfV1w221+UC2Dl2yJIZ1TynzYypkveLzc6NtG4jnX3mRJT6
vuEZW38LwSeS3Ut5IaGmZ8uugNKqHqNAcpTNYVbSHkh1End7DwBRTmVcWiz5oPN0va2f0xvgk0EA
YWUrhXE4Ht69RJbrQud90FGpiOO4XVTIFEC3y/n85pZkP0QPtPMd+G/UinKRu7zy7X/AdvtO+oiB
oxqPYJSxeuRu7vSsTUrwAQEl5DO3SbIYiaMSwrML6MrXOa9yyTgUiyjt1XHah1U0jzMbvTI/8jBf
LMA01n+Q7lp597PUyzWEJkTgB/4LfxPc/L0XxArzxO+mF+PhsaB+NnmEXD6hdYEA6B2QPS7lyLFI
K2vWz6fIv2cI6Q3Hv7ca7husqygurql6cINtHlqjT7d6z8g79qb35NGoCNWiYFAGWnZCF8F9UKdm
jPvmudlu3rCH73YVtSGqgwSrZKPJIb0c/YxPJpRpqKgC/hN4fgorJ84MmLTqHEC7b2xYlivPlMYj
vLnx/ZNeUv3P6WcrWQS20zKXVLD8rD0MVwoViNERwrhbMZatCWCN281G4Xx+qxbZqduEYTai5jRI
QB5AxXOW53FibAUCFILffW72Mz2FtM4Ldk4D88Voo/2prAcNO6Obwd61ndaXJMAtOs54JPXs8UpF
QetHCS9nZtBPkCsshaozcrEsPJ//M99Kj9LJiNszhUgFYdDF8zaV4eMt02DcCHJTSU32D/A28rdC
iVAG8kEcv05KSH2fH23UqjRrDFSO0E93DA6YCw9bm3nb0IV1y2rSzB8/AuV3F22kiDh6+82YAQW6
ZF9vfNhg5DlL7avuAu9HurgmFOiSoEfymHnDKWpFddV85pUFRRIoYEM2Eh5tzJqj3K7RgUwk6meH
flPi/3P1QDzOn8e+jlDra38cC18DylYz50e83c2ZJBh73eu5KkNG6u8mn5TA+XXFtJW1+QOE7/HH
DKDJD3bJLle6vMe6SSO4RYnpngG9Vvzd4vhuJFk3Z7Od/QzESuKcue4en7l8sEUYVC3nqmN6+u2L
pAh0mAUTuJjGY2hLNWTXbZrMDtOMz2YM6Xw/pyF9vJPpiVY+Qq2qMnw0Ww5bzxB9Ot+LFSVfszyx
0yCRKLl3YLwMZZUYUZWeBIPJMnvSKqk7HzY2rcGRgH8GPw232goksN5bD16QuBTDECfEDiSa9vA4
bXMT+k0M2F0nKQEBn0z1bhpNfgoxYWe4Hf/h8nXpNvSAX9rx5yU5X495p/CMrd3p0xLINRVaiOX4
XAAWTZAmPrue8F2an1GFD8HrJ6C49H9gbgl2tieRNHHnbg/ZhVa0c651fDItaAVeTgChQ05H9C2Q
tTAuXzXdTInR9zmpHgrbBlQ4UdE7nLl8DQNY6r0xSGTSITge2BY8ZnkJyhq8+vw3wvcI1NkoS4sA
85FdZM1YAUWPakGAPIFu4Y3EqxIz9QhQIQCUgX+dPeAGAT+iAfGzuNSp929wJdfHz4ILBdWSyg2v
PrfBIyDGUKUAPGWxx0/xVH3F4LVPBGvHpCwXFmttJc+l9m2gp+0Iri6Yk5dKEZl4T65gtVleY8so
DzaaXE4zuGPUFBeKhfd0LrW//EK3k7Vhz7fhBBH2OVMbN1sipwJEZcufwPN7CjuK/N5rCNy2KAO5
9sVdrluqwCdKWTFkScDi2Z9iAnZd6JtO+jLNimwxxge8qw2Qt80RzcymE899HS+8PH3gHY+jM6HA
Lrln3jU4VQtAA00YYTcyQ8rPjV5qAbPGqneeyjMBs+JqKfc9hZc3EZBVmk2A2Fw3YJUUaM39fd+0
0QEACIMqWV3w6ARmaIDcgw28XnrkvIcL1gEKxQu77CLgDDHVLyHx4fQN+DXRwWbuQiRwR4vCf99d
0qNfxLCjI7moeU874p8Y5AwpXJTOhqL4QGA5j+ZIELdl9KYjHe3ScbULA7PjG3h5ml8piX+vGx4S
nOn02yPzGDWrOUvP6SkknW5q9VaQTOX57vIN/BAbLOTRjQTeMq0ivoPByGoIwcM0BkoXg6Scpctm
tsij7R27UBB1QG7eqNDDim3rRGosiOM60SLdrmfMlwGtx8cfyAXPJHCNB7fe9LeCi/jYmQ/y2Iqk
/jOlDP8F0CZpCxN+zpKxGRtAsSW1sIuNcax6oy+ZclEx5Kg8i8brJuz+ZRbY9Rz6fgbgtYwakjxD
+qivvuW74crRRWSkYvQPpynEmw6yZKOAh7FYLRmgOTLNb1x131hkCex8MmSZHHptVMyjS/8dhFoJ
zAY9e366Qi41MtbXACq65XxQdUcAjklJ7Turk7yaN//ydwymO1jzhQOE31rBFCLPsERAjwLYl75E
D9BVv2o84/xvX7nMIzPChMjcFungmDQA3xtpTWBhiLJHMwUMilkVEPEJINaRkZGO+cVi+NFFIBRU
yiwW+XR/mdM3nQevY+Y6txjn1dwRvSf8RR0NQLEVh1AFVcZIa1UOGtYUHm23jgKTuuiTjs6MtSaR
YG10koBfHne8rw3I9lgwKMPXrjGFcZ10Fi7y2vBgz2GS/7qFpQHGx4I3vou654fxaBWKxt+z8R9E
NpcykctqYSw5kliOE730vdmcainjnhlz2A1lb8bbw0Idqw5etyCAZYPPLchpmCdWNtSAqnqukF/Q
lltOS+nVLV/l1QWhOUUCGO+dW9f4stjxzNxI0azZj+tfbRior4wuA/vs6vfleISTdExi0Tag/HU6
K4ZmBgTzgeNoX4j551rUyk9FwqxWu/9Xo9MBnDMB0AUW7Ru7bnfEU64ejNz/P6CQNTETNoQGb+YW
8dfI6oniIgHZ/qb8y44CEJnkXPtPd9bLMSfI29lRNkXLV0UhbuJz88bI9Z0WoUdhMtZWpaPOLmhR
s6Tz9gB+TYAKy/DWokrewTkqEvPSJrxcdZf2w+umUip5OF58smJ7i+rnSigDZPMGE4rG4cJlXCx0
TLSkPL901lVe9SBYI10/cUNPgiBfBy3+Z7kND567DdsqVOVlnl4xnD+Z3EMRmlQTR6D1cNye7CT6
v5JLJ3AxHQT2DwVtSiDHjB0xBIBX+/AMNkzqG4yRIkhzJvAe4Tk27Me7Yw66M3ZEEo5yhvX9kQWK
Gf594sAPBmE/OpKB/Vw5vCtXRbl/7iobjzhdhbvXmaL5M5LQ0YQZr37lUzgWl4T/Ys8JtR9KCoes
LcsDANIVDnYrSJjFUrk2VmB4sfxUt1C1Guq/gj2UN/St884cqnHR8pHs3TiuWcOXO4mW03DnXShS
NeZGASd9PjJ6WtLw6Qy8EN5XQ0cq6Eqibwzxni8EZKuRpN46GywzsG2JIx2RQJk0fwOa4Ft8mdYT
8V6AaOoyA5juXl5xdXRNZ7ncni8CY4yqFOM/bk7yM3vmwJx08d5I2oW2rOkef+7Pcidf10YguZlz
O8wRaT2rMfOwbtUybsh1U0uGdKIlHwHTjdGtlgdfMVrjQvJNuSJmqc38jFTmf0swjGif/nqNo3ll
GoRL5MYGSggVoOSC6ouE4vtK0yR9MY/6oiZ+zM+7duxyJU3V7EnvUsqh+LWKbhgF+0RS3C2/0Aj4
PT8kWcqUAzCiTOe93kYMGDfHaoddW9etBDXFbrhnmYSiy+GBkB1L98QfC5N7YWzsAtMEgiqOdZM6
tkIgi+ddY1f9Ny4KVPtgIf27YvvtLDp4YHQzIU3ovynFqE2iLlCa6dz+mAFxmm9h8s2k0WmYk709
mUkhI40hgf24saghNPhKX1iTokpG6oqWoscMKipXKwl3AdUpQei6f5i62L8GNogZME60V8RKqhnK
P5oGdGIRxe3Q37bwp5SGADfmMdLTO2iyVIih/YviHsNU5sB/UzQ8ozXOW1ghgOXYB03pVNkOeKN3
r7ky+TByFZZMlyNL4HHen43SyAiD3vC1QmMkn3MndN9bG783XR+eTcGyVimEgGt8o/Nehx2yTqk/
Ww/v+c+dDlpzMqFl5z61rritf3on5zC9jODKMR+/fMwgkec/HS503uttY92e3GYptZoZwRWyiSc3
KGJoq3+x4ooWo/iLzBvY7bBQFcyvyp5DKnH+qSurg/7gTeAzdVexOaIf0G68ta4H52Fw11qtWVnn
qdb7djxr44r1z1p/n3QsRDwaFnXFY3+eOQGqngYqGXrGWivXlk0a0G8O/iqeqOtOUhsYp3PUs8d6
0oiI9UQ6O40mwzVTtyt8Y+TOE/S6+UrF1EqyTsQ0c2iJ9iJVYBmAkbVfT7sGUd/7GoHM1ezSppHD
wslnrEjmEcY1967NGWKPpDGU1gDi4WNEEeLfrc04I5DDNU0ESvnaMdMVltMMnIo5VI8drWaCxlqt
wPW/kEc2VQdVU7sROEFTOnI+0sHwuioqnZSVmG9jGzPmy9/QuooNTwn4lL5xLyYayTRut8zFnXzj
k/rqF8Nx7hpnkf+etaoBxdNOVYCMvTuJyt3EscKQE5AIJk3B0zM4ntbzSWULeYJnpAvCCHh5P0ar
EvX6hWAXFqLE0HvhnKypPAOUJduFIlRNsUgtND3wrx6EUdrZyNbJjSOCDG8jTUfmg9OPQslviN71
OLAQwQTFwm9M0a/3RKWQLJeI7goaxF6gJ2fnvOahSnpSPhiutoU/tw4ybtFBO58MLoqe0L6J1Mi+
lUreEnAJLJsMhWtPTagdb/tp3CeIRQDBSGNOkVheR85U3tzlo6uxooLlzAIf7TLElpdbiUVNNSqr
kwotsT+cTRHAWIKd/hPIs9jiJo5Dfvk61mQTQMixcpQCRQWp6vrL7pRKjJifsq6GzG8vqkVRKn2d
gxn3GhTgqVmHI834uce3E5YoBBmtgjpU3GQ8sZMawVowykmfh9BSrQjzVJT1XRiXMNSwTsYGKunm
gFp8j9oOJOtBoOSyUNubksdGdnqxUWG1VH1EJpuUmBUzEX7vSQSVYNZ38ik5NWXePDOfdBo4FQB+
le6x0/YnRPZfwAkpOQBmK9Za68XhTseJtfQMfmiYkNR9/WXk9W6FZ5S28mgOMWlPsBrc5dpdPByd
jLZ3fX7z7NDRSH5lJ66cq2Pruqbx3ET21C9iCtzbyBTKcxSc2yxgB61ecHyQKlhfHsGaiGJycz1b
WrxCtkG+pyhSqxhy1smLpcwwL8UCzQwkpE07poEGes8xJ35r24zd0SDufuqI1vB407jfBEGorLdp
XVuhR5ET3V4tDpp/MnZJfOgSFXxw9HaskOk9KigrjNSjtbS+WbjfxDTgijxV36wElCUJEg0bf8LU
E0iBCXUXwWh0fTEPoc1y/014Ta/o98yk727LsfIZ1VJzglhd53YP6CcJZ47JksTOOBcEnT6twL/l
0bpGWVXY9XZKxVKjX2Ngnz757LafYl3T0bB405VvJRQkWbobO1KPDT49GVUIezDMZbgZvfx63C9M
BUyWe6RDk7qyQFso31OmW+d250Tn/sSjgtCSNYIx+3suzms8Kk9Z/TU8uWnCsc04DRedpf2FSivk
A41L1Y9i6YTJsJUn05vgviF0pAoL4E4YlKAXGBysL+i1MDSDg2dExixJh2o4U+zOvxmTw7gYO5Vu
+w57Yqva6ADWpUeBLM0fDmun4G+/YYZ0cbg2KSp5otMC6hzeyBbB/8Sozgz/xFRMdIN38dmbjJFK
fBjJd3qjJZzqNucu8z919C8NElf3UQ9q7iUrdhbuX+1iXZkjuCeg6UT2j7Zv4rEex8QVpQ4qFn4s
un+gB2fBcWwTbWi68uJGGYeJ5rEMSZhP/s6Lkzp+l3N8VkAzeYfNPr/WnW+PHh160tqzwyt2QGtF
a9i8zK6ylrM35L1DQ5k6zVnbUWG6/zlONsn1Lzt6p203m3GEtRJsjaiPZkhwZsCdkVaoAMx0/vL+
oJWA5kH1vnuy1jCo9Ygwv+pcxSJpDi2iHtinHwvmup3b/dWR+jbXoUMLb76V4BopkQREOTPI2zzo
mmLtTgqweYG7GjEsZ+MRbfl1bq84fBhFECDT/jKZA0j9jvHvqHwgU2bhpDP9bo3AP3350vgHET+H
0z+xY6wdhlKA/Kj1FQ9oWB+A8iGZ5uePJHQU/Qh7YnBj96CuyCc0tF4AVPKwEp7l3Sc0Euc06Qj/
z+3L5ors0SLRjPv11R+KYSjQ3zMy5vKqH5tKj7KpjmqkaUJildHo8AC72+VwZrKkn57uojx2AdXY
Oa67Gdu3GT+ZLc5JePiBn+dBdOqGz2ZDn/Corz2Y6SD7LX/3VskEtn+vbiWx6A4AgKD9mmwVKgyv
FfYu8HpxXzZZL7mIELSEE92sBxqBvEVBX8FSNCBqoRCZMqQ8XSmFTroW4KyLU2STxk/C+8SQoYOS
8BHmSv8hp27N6QRa04H5UqQsUbKa77h5bVlYNGyNhg/sofZbmlamXcpX4lhUEfBDaW10h5Gi/DaX
uEjrGHOEBKUGUsojYczLccGbokXNSRbyxG+YX20yckjYIvz+KUBDzoA1fAgZigY9EL53idvt/bQS
w38nquPYAdw1JrT80pxz8nGpPf4h8lqgCxapHU0ylAewU2S2Vid+/0zuusTweN4D+tKi5ycCx9k1
HsjDiHFqZwoRh7d33GpAJ2Pko3HZJ7wAwBnUYu+YCRjhqv/1tUImsvF+EPKz8hQXelfM3bkGwEtS
qAU+t2MqAMZXIF+i1aSdOyeapZx+rLxCZjt6CtZ2hdCVBcWqq2XTvlQZhZDYvvyEEKvVAUrl5LTf
+2vheWjiRiH6s9DsorFUZoP4qNLzT+hIsGv5Dv2ufFifF28B6aCIC2+VXWZgTNh+/8bXHXgZq9/R
wX0BXF0++BGdty+cdS5LPp9uspawf47xBRFFrZsSYZacrFnGJe9dRkQJ9qJj5PhS049SBiz/eIKv
atg8KGjVt0M4qT3iPzRvUdzZAa0lZ2BroOHeEjQNKR8Aac7XubKkWUeeFepmLStnI4PV9DrdxcNS
r1i3JgoiL1Prwems+1CuipO9a8XWYINO773n2Njt/xfUDkHBMmxISWMqqelq+b+bAoIcJrDAvf/J
QDt4lvX0aWWDc+JU2S+G/8pOj07iBrMagRqdALGeaMlAddd9BE4+YXwA8dgJyOW5BSOXOPBACNOk
w+gyxbAy8kx+EJ/EbRwc41Q1UZErgIo2T3CalYwMlNMf81ER/PRV8AJbMIumSqGq9xp8oYD6neNW
TePhGbAXtTjGEUcexj2srAxeFGiDeQ0KaKA+7Q7l3dU60oY34RgUSedIUWW5siNv3w7w5d/7AMgQ
wZK/qtcCfu7qFdCk/psjLzH1pgzV1O22zqRYJB9e5ppM/exczXF8YbA6QhuMAwqaPM1ph6shTNjb
D80rmbC9HgsQrtClMWS0Ntqct08Izml8PWgUYhQCezsf9J6WoIUUOZGoqdhwiad3OKCEpTPoafWC
5DviFfmgnhIHsQmO8PO5ZcAe0N8pz2D5x+c3+fQCEwrHrq0TOBT3DBWjiKAOFuBO8sSY+h1dSLrG
W6RMkIMSNGDQFUibhsHVUFlZksGFPPpXKwOblXpHkQXm62VTBQfARa75JSm/71kB43bYH7FgUFc/
m5+ashkge+UFOclNP/CcafE7gEjTtFBiyg1G7f2aw1deCL0jJsBydJeCvyhuI+0tPdA54Coqn+AA
vjjhq18qoRhM9kW/SulhzzZdaNY46fsdJuWVp0lXyz3WFrblHj2sRasM4kV7bnOyjFIFjnem1pSk
3/fXd0LFHF7+IlwnptCz/ETDCKcl3NIGrDmOnr+zOEZmH1/rsWnkTq6UBrweBgWqKLWz54nOSlk1
oP/lgVlZp1udqtIhydkRm27U06/zP6Kl0e7yiDIZDI1o3RQ1UpHw0ehtrtHuzrMGXmDwjZK54Tkg
yW0+s5L5ZbTDR+qGrXw4awUdLslxXSffvzR8XLyZ8/f0JCWvF2UmwVbMn/1OBOhWSEKMbnNsL7eP
ah6v9NwGYoKgM05xxzvqcMFnfD7LRYeoT3b0LpWW0/pB3PoODMt1GHX2Sxt9aCmKjo1VB7Cy7BUk
H1RiNwprssuBBxq44QdkSpR8OC8Ks0pe+vRnnfjDhXkAwYbouzfkkT4MJ9RtRn8UNHQNwgCbXdHC
BsshICPFM7xG1Fi9jiSYr1r6mVuO8NmH9k68r1SBYl+H46VgGvgF2QBDOscft4C9zJKMyxNEOCyN
wt55eOshrsQBwLx59h6IohvJASHOwPZAz6RS+u1K5cS2euO18G4NkQumMQCoFJ06tSLdO0YbXvS0
A1PaNV0jLy1i3mOd4x4a19vFDBUm+PkCNgPLsMzR2uIl44Ahjc6SlJlM7LQ91NucgTXq9Q7d3CEp
BxEgzTwwrF/LG1LYD3RiQrmF0lEWUWd4sV7uhKlHZZ50PPwcgJWgFfSNsecORrl4hZzAbGfLzCdD
V9lgwoFMUrDosiaBCVxGlkU/MmYhxjyzWXbbBNve9rbB0cB4oV+ueoT23oy0CoD3VXZrPNsQUpfO
8ZDlFgtUakcfbOtCUEodb/9OZJSn61W5ZNkzFLlLhfzH4ptB0CSJzqTV6+exWZxwqoKt+LZCklTZ
nhWWa++hgJvOH+hktuU3hSw4g81NsEAs+4E/Wo8UiLx8F8nCaN9dEY3bmLUvofx201n4/2RIvJM5
LX5YLK75qgljxvcQE9vohhYzlx41O6lyPTpOM7VOAy7N1Q9n+Eopm9y+uj+NM0hB5qdYCGLWCwA7
9w0UrYUgOO3vBFPleZUesNlfcu7Ru+soDXUvDNVSdViBaddpCg/3od3kIAo2BAd4Dmx7YSXUdGKR
5hqvqMzurjpm2ku45fhU5AJKi3e0zQQ8a4rZmPzMbA9wmndpZRWw4X8RhLSZI2v6OBJyrzCzesBF
7jXZXefm+FV5xd7636GzdsRttC8u3EJ4vP2wlARi3migpoqo9zB+a48TDKZYHFz8LbIi01NIcG98
UGsj7UCmMV6CqSZtDYk5E/lzhJtIjlG8IhgOl+qw9jeM0JWzbOFcEOfDXuQZBVChdFrl0ELbLuk0
17MMBIGTKz/XDR8ANfUdVCARBNiHBm+vNAyHK2fBqi8IJYPbRHJl4FmWX0qlwO4gpbKpgD/r14F4
842RZbpTgwk4Wd53y6LV/Zmnr48e6rFmxe3EaugG0BxALub+8V0e0fHCfX/pUb5etCNzZK13pM1n
WJljdMpz62/VUxwC/xxZeaceJ5OLHeJ0FMPOkipX5Eaonj0wRnXdvXKtwUHvTyWgskr2Sm4Wl3kW
yIf5QOOx8ixHQRHhajcUq9+NXBJmQDVs5PQUiU6RPkcOQhPDNDKiSvX45iYVj31xIj61cE8DJqYc
bWu4qrVSo2+bpG0C7R6KXPe2RCnR2WUZ6PgSM4SmR4Ny7zeVcMzxGUqxvqbKkkubTlOHCOUiwzrg
NisQ9Et0NKBdaeUsJ36vRQSv0zBQC4ek//sHeNDFd6VfUBrGLuxh2pHvGA0F6+01Yj12WQj/EHXi
B+jybc+mvWbB2VpGQfQ8diGe8qZV9yse1dkMH+RiMIJbqAWEb36gLRhU3Lrckg9MVfixgoUHaZRT
hkuLzrUtq4HGgZcjwoE4gTVYJs6NqNNignUy/kWoJEOE8Mo3Bv7MS+zUlZiH4COZoeZKiNJUQwht
bxPjxQ9U94o6nqdnE2Xab7DGTUOs+vfYorOrqMDNHZwp8aA/zTm5kxDCyq8xGCoiBjP2PZb1HwUN
cVmGQ3NSUW5h9gwL5SO+VW/QhqXaAWrvrxoxf2GBkEhshfUUePcCIQOkaZ0H/I3ZxuhGDe04GpAX
VQG4Nfv5IzEFAZCs6+mWKFbsXg1QR2FPHzc0FFahyavy5M4XXrwatb6avDjdgOBjkm+yGIZMQlFD
RKT3fq1vugn8/22R+dN3WEFM6NopyC7CiNrXAQAc2zGBBq2OL24oFh24+SuvWRGReVcp6WkyBJ7S
Lams9W+EzqvjwmvdcFASnZ35zKGV7EBzZsp13wciprrJAT9mDKjnc/EnrXR/OL9Sn1NXCx2sajyI
913/mQCvfgSB4INZcqtHnZ8DHGLsLLTHWeIJn1WLdmB0MjV6rGurVMOEOjxFHshgYw0vzBGBcCyP
bCli/o3A2rki6fqExTz7aS+sum1UDerkksrUY1OJGmTDUDJg+0NdT2oElEWkkK/YNlPSfK4J1S8j
vDKVTvwyz+b19ZPNFgiQPkf08IWwQAx/Wvzq0dVjW79aVQwxd5KGNfIKkvKuP2DZjm8jjxvoJvcf
PwTz7y14L1qbkV4ZQIgRPqfqptm1MWMjZvHXwAUhcKAdeKc3mEQSzP1wQTYsR3k+Ujc3StKgMOxP
qqegwH5ANJfsZxFkxSo9d86kw9oLH/TCSw3BM8peHFSzPHXfc13HrfPCklnOvR4SnDUVeFBNUD+q
Ld4Aw64nhyJRaQErg3iK+/EY2lylL0zxehNn2VzVXvbjFQY6HrYCF8iVrboSfmn+hks4ejd190b3
WgeMTBhh1i099JnOTM6akd7yn1+iNmKeT2fl9LbjswonC1eaPyDOBvzCbFHesvnnr6hPoeFjjJlZ
DvblNt0JgoFk4vuwXlaknmkitH7gdbXaQnKIpxYVsHmGrlt/4bjMPZtQxmBDvKS4XTtzHvfmHtg7
23xd9d7FAqn9Crl9U8LsFNcHOKkZqpj96tyht6H83clKEtGo1IJsD2MThz2GzMs/Uo+gjPUA1jut
JpK9D1pmgTQVdpHs0CTt1vPHx0dWPFJZpJ23dbFLSyVcZPN2e815sMQG6v1I9MDvoGAl6V6UphAG
Z9os6fib5nK01psrxcFUmJo/CR3ztWb5ZaNlEz+qOrv+hnATe25qeFxSCkhEfVDh3EMFuMho+KfX
vu5QC+F8AhFRT3VjEkIUX+JdNsAMGH6ENZNVVx0z0DZc6R2KEZOZhkO4Lvx7B+h4DXhYeZ0F0LBl
v/31sQRihpYeEpwcyoyAF1udsB3rUM2cUkP7LPbVXB0qVL56/hk++b3sEuXQQ6Vr1PNaEvofm0l1
yN1uCPU2AVMQX/ndkxFn8vUkoHCiDZwidNL/JRTHKQV2lKdTEukACvCf+Md8phz9/Tmy/iG3k6vW
QStHH7zklFmhFgMKyMaJNkZgA/RP56WMwYnqz2Zyn6qNJ7VQvvxf9cKaqMdt+laPPeXyMZyROr/9
W5eqvwQQhPHvn/mbzALWWnJhYFNPXTJVbE9MrP6Fm0v+NCuNIMlH6JxHYHh5iCHttFQMK6Z+CXFs
lJ5xqBEcVTR4Rle+2NZVMLLXP2yr/dkXsP/6rK8x5vcFuGF3FKrEsCwOcaDowYrCfwI0nlQlSdTv
q6wZ0PJ48i+WE5SEOpGPyzq4g2fHqqp+7QcIZM9Bki+4ASPkKzmH3ApXMB5OI9d7W4xL639AAyTn
+KQhR4AW6MnG43rtSj2DLYkUt/0kITlWrgvSCxjx1osdy28O8lLlWqvPcJQH6Kc1EEmHXTvZ/po+
+YKQes3U2exe8vXZWTi944Tt3uUiWHAeJAeH3SEX7VCqmg4i7mIKyBpKwdoPoReLb/JzUxEhr2cK
M4o95zjd4UTlkhXnk69uDQxEtwaNT20PlsExYZ2mjbKN8H5YLtD+hcjzfCdnptpaJkQJctj6cz7g
2oe77Am5D9J4UJXpwuMSGf2QEglXgdu7vcPEALRxmRwt/y2jEt0FKHxL3m6fpOsubh12WF7itsEw
vJFcZhYxu6RBADJsDuX6dqpTngE0lFV13kcyfzw7AZ3EMjbzpSMQ/KE5icSnFOcwYcwvTridnXrJ
vzqvmIUO7uXv0IhHIQ/ZoTnH3HfuRuzVtKY+c/8QuBcJ1EfNlE/cBfmVk5+JbP5vr7XqEwKgS8+U
fOI6WlKVWcC6CiBYKCNH0BVQPLE4b4SWqnsIwDpZQnLHi7x8eYmGxhlosXbEjvVRnUuVQrSLjmzx
Ti5PrVG/0bX3LhIbev0yxaWpmKZ7NhxQL/2pfl4NU+ROkmeYW9QRhXJ1IjVLkAPZZzW/I9ibe3ny
tcK0KGex724/gOa1rhaT4DtDXJx5VYZUOmmIpoBXtntLtWRrYcSDjjoui8zcS2IvU+GW88b1VxhD
a0OdPSvCkUEnuj+ytvdzkL6e5jqyUg1T3CTZQWMf22Cfimh70kCoQauzYLVzMEpAuhA4CD5cQ4w5
Rpy+FKxrTPZxTDMz8B2a2iBxfsMSfzb2bnQcXPQ//IT9gi0tHZgU4B4bCB/bUatet+kXpgaBkdKM
quPC1u1jtXgPZ1yU3wCKMZZFclim63cIcavWUSwcSSxipLPotste4+QlipXyabBngaJCRWYw5CaK
ADBPS6iVJPCdyLxs48JPXe3Rxfxy7STigAFHIWf56IkAs4uyjj8UMQlo/ATw2jY8c4Pl4bDoZxye
mOx4SmPGwsxHy4rjyihsUO7XDpI2siadi/tUbOjXghCho9Z/m3WLCjDE2jtZJ3f7E5Ww0uEdfydw
tIgbOR2CfVcE7FIxz2v6vDPyxWxMpn31Qu78TFz4+tIQbO6bo9cup+Z1ddhzPA2RXNfFL2KUwOT/
eoKjHL2dMEz4N7yACfElWzJxfni51uz34eTyEd/f5ue0nulxPuJ8g74DTzs1med3TneNuX97v0iY
80x1adcxUhdWLjLf9oabikMV/7eEVjP+HP+ugipq20MvL685k5+kgHykk6O7zb3qyKc6mtXeGIHO
U7Qw/SqkIPP4ZYUGjwIr4OcjLRBlwNBG8zFDpvux0WpIpvV0jFmSaiiZNLNQLquZe4cXumf7C8/7
QAwybDpvPQbWgHYdDWDgfB5Smkxmri+8cUJ9lPxWRsmh8o/30cwMel7qavfEJ0OI1jpNpJGJyam6
6fll+WsJUkrw3+VPxgC6MShmrit49uYXGEa9y/+EuG2oj7OySUHt3/DmmdyJtowCtYmTsXohPqD4
NVebRjV/WZoCS2w7F9QQ8Z7WEVC6O2iBetl30Rl3nQxg7cPRRNPr9xiEW6WjPjGHNSRIKMGPQoTu
Gj9h7N/7B2wnnWC8lzYtZkgHHRhYI0zg1oKxHbU5s8xfFtmitTMCBxBhok8nPfvriRbBzdt3mnYz
h6LEin5YIIktXZ1E1WkJC/TRnW7oD4Q3icEAUt+cZwcD72af0g+k6cDX8nOH9qVenEFpToBlhGZP
ucsSPanZXazLc9QSOm5a0KrTUE8/TwAqWDfZ3ccxg/KfgMZAxZKNvqWPqMOYEIOaWs6yrRmjQDls
DNZgqa66xQg9nt6RoeSBPAkOchGftV6s5q7tR4qSHtjnUn3+30FyGlYl0Bho9L0SNX2uGbA671+R
EyhCcnZM6OjXhlNvFFPmYBKk3UClNdB6Nmh8DiGtlVCTmuHufcwhGF0GzTWDlQAGJYQbSHnZGTu7
RkO4VN6SIgQiZ5esNUefNdnV3eYJXzhRXqqRHivIiCB79FQCRkxOsXhL8WMvRHHhmN8VETyb6lF/
L/yUxCt7teklX424cjbUjsSNGVlBsAeOLTcni4LppOdkdKsza8b1drf2MQfS1rnqLKk7DmoJU/eB
L6ZCEd4eDBiQ6z7v7OvTtHZGRY44bOCTwg7epmai6kS+/YscL8YLlg75iDguJZA0OLw18IioMeYt
ZPENzQL2IqYhSrEHDkc13nEQc/xXhkH08UMXAkPHV5JBSXtlUHr3YHuCN7U6w75uuHBa0CXBHO6+
rpSFOU7d8lKcQZTnwG0FbQ9+ARh7ftOxlFqYKd3NvVVfOBIDjm47Rh4XAllPBTqw5w1QgJDWWTkM
RQTyGe7W3cpX2fvgBKl1UFDfbqNCr3V0+cPEec+p9F7xAT7IsrUtOgN0CUUu4Gmyf4zWhRhgTrEw
maeg6j+FD3W92g9/bl+o55aDgj+F8d0Ir5sRZlqHKooB4P5pJA2R/PFA6u7xODLa2tKT2kS+32zP
P8QNFdZSedIMgfJG33J3fELGN0kPZGdafzxrICfTm6KOR/JNA9JcqDLyn4a8JATFkxDea2IHRoQg
6iTVCviou+7PpM9EeTqJ6jlfGauRQyBgDqTJmULPFOJh13XG2adt9bgfrJhZQTXjHcD8sJmaWhoa
6o4hXi+QDLKRRKEwIFZZHAzA8PpNSbKIokd38+HDDRW0T8aiCC/nn2MQjFlfnfBa+Aq8kXQ/MWu4
G5Lm1u2XzYCF6E7W1xNjq601ZGtIU5iMSQPf+iJelCFncruwOwLjpl6Y+Sx5aILstauTNxt1h6ID
A4pddM8KsYyC222ffHm1Q4xk4W4mboMHVKrIS14wsFwjaiA2HkuUOXJDfjYO2rYyXLCnpD1s7U9b
jZllZDqPePb5eEITnx+x2BHxEII9yksc45jHptfeiSZ9dcayyOEysYF97ZHA9YQsaVKb5CtDJIrx
loLFNXmFto6tdARGOLBAASBFs8HM5DU+UUyQe3QuqFxK+ZermUlgWT5wXSlhWUPQhVR7BesSHiCU
mNdXi7BHJcJIdhbvlyLg3BWDS5PIwP/7t8VPQLQBqDwdNWATNZd8UFV2zTDb0Z/T5a3YLd5xJP4M
g8ixW3KI5L6a7o8Wm6RiSq+UUVNLZPJkyiJUQ3d12wlyqrl5dmdFXXZR2PsHUDYicKVp5LccHUgJ
4HV9uIZspMAUcyQDC2hvChigMcSflRr2ZZnUqnk3of8HSA8IvYTGf/N8yCMtC5SVW2QESXsvDsi3
+XAkW0fWqxfmRlLoNsq4dBf0LmPDvymp0NLalsgMA/nt8CTw4DMrccV8xbtY/ulVM/K0fLwIhGjI
9x/wT63lyC5B4D28LRtYdk7pLpWW0Px/kH07/UGPanR2Q6RSF6xvjimxF/XvlDnsvgjdNoidmOhO
Bf/SbWQZhFRTp29zVJkLoLDI5e6tOSTmbsHOpoPney/ZwbhuD1taccUbGGhemIfx08z9dFqqj3K7
xq9u6N3jkpLVt7KYOPDreg3rWjSkXTIwIP7F2bXvlYGhTcqoZvYtLPelMTxvyYeVAyV4sR21mzAd
Ln85nD1mZKjhFSluxPr5tr6T4IDq+454mWzmP+tZkciFU/X12v/3xinP1zKWRnF0mioPVoPdVg+p
fAUTcPlfLgTt/vFPZqKiWbbOrndmK/o32Hv3RXU0Yaq1m4S7O8v74ty81TAxsSQOBa6yKfi9myf7
YF4LhNLYJ1xpTLn3hOlVCSGWtQZ0Y+7vrIh9uonm5dLzGEaSw+pMZVnzV8aTjB4mWu7Zx8yPbf1r
ZzKg6rGe8Hw0bJGRL32HJqsF3XWPhT3ELJShzaHGPuoDwMchW/0SJe7Kbj4UCdKVFYblkJMQF4px
I9PJtH9OyRTX7z9z4bRSxi4qDCfhetVYN+1U8nluL7PEr35ynSQXQNqAo/TG8RPtsxSo0dPLrA4m
WzYHZXqM7dRzvzrHn8BFBt98HG2yMGspYk0XaD8DQWObAd6XlwBQOm7wNGDP4Ajcv/TYJam1KXhP
Fgz2n3nzQMEwoeytuxd4k6xHi4keWWElUr3mcuasMrcE6jCVdaupKeBkFSlNsmAqM7O1O3xqIQq5
b4cPwyZxdOHlX/VO38+HT80Q3s984YWQIaVtPK97+6qC9BXrnRWRjq8J4bVP/AIfIp17q8XKfxP2
G8TP3Wju8X5DRmOVVy16PpXKxPJw1CMtCvah4Ozvi5TT/2Dd5FUGrM5EbjOcrU4vpFcRBABECevs
VfTZARkj1xCAJvP2BPlMcAVKlidwpQrTshFcfV8drFXFwsGA6yqH5bHkcVdVuQFazaFutwxbHBD+
sizNdh87tNY+zkYd7imf9dCdZayZunVdUFoo9FWEj4GC5SoHM3g7dKU0MIrftRPDupjcPahBAV02
o+mn5voXorPESqfkcX12DJuMOcxMFI7sflS7s6A1SqqnRUWIT592hPdEOntQthqfabVGjIdmPkyP
+Y6UTDniYqxri5Zib3c+F+4tJEYpuQay/w583SzDsaUbhVPbKZaypeQCKnyRS+la7RQaTyuO5jE7
mS7uSNNla/ECdeeu/D/NV8s8/+GEbXAaZid1wByh3wrZOTHp3af8sgb9Ca/3e+2pgji4+867Jf8R
RrMtUzfgoUaVQ3jZ5z4isSTA5+i7bv73wLpagJGuvu6V73HpB+95tlJAJwv4mTfPVlJOfbXm/lxS
ITYe5/7W+Ae74xfdh5/Jp8PlVxH6icd04asSfooA6vQRlZ4U0T9YMw0V8s3zs5T/HoOQ9F6PgYJv
VeF7B/qCmv+hz3yOtIuIZtkuxapwREovjR0WElj/r7lOOjRYBqHcNT3dL8tjSWn1j2+CKS9jYHjJ
uUmsqeYe9aWgXOOqrRXbotWkqa47QzbsqqfJoKWpGqdKhriLPfPgV25TtyazdLZPR82xge/AMue1
QTRO3w56dLZX4XDdkcSCJRP0W3vG9nWDhIoHiauK5VNZHYk/aM9GJBpLafX9NtM7Qf+U2QE79g0P
uN8asjOsFIxOumg0itxBb81tUhTxnaN+HzBSA/pf6LHWsQkQo8xmj67t4wKR0Fy+Uk040F0JppR7
HBHUVlHaCnJCxg5S3GphVPlSWiqYvjf79PVH904nNUPdJPWFuPmwLXsf2nmtl4t8nJIAGHJ89N4I
XXwPehHSii4zYQgbc3JURZFYFNTQcLObsyQ0wNCKMXdGR0u4B/kegRRDoGCbU+0/EbaCjaAnahtz
U1iM7uwWfD4e1W3+JE0cvECE7oRoYc7GfknXd13pRm2HHrnEAfwiG7Y97C+ayQZUa2bXPf84GanY
W0xmuP6Czy1UFsxAt2SVKOgbKFK+LLPvkE1M8omksW0hIuDefjWPQWPX0/6Rak66Mu+1emzTCfww
pnSQ+6+AWxNgd+TVUXx9MfKsrO0wHCNN++zBkPuOWi+84wCP54SgQ2ESxPhrakYuESnDJpRlA1zg
CL5byXX95FWK9PUS4Q+L31PDTBSA6X44oFUdFPztlGSQSqRk1KG+Oant8ezUDSrpAKioCQXPNOZR
UFevoi0/ecx998urpCPz/Vl1OiHR5R9Ou3RbIiq8HUW3D3+dyqnbsUQ//cn4WHfcEtVDsDYWgWFz
ru/1/aNJlZUafrtRPDENrUtl1cUU1qDdsztotXvJC2VZenbi/Q6bp+nrZvF1XjDXmmf3R/aTd1zm
aIwqWziEkZX3GkXqIRN0MgFC2aSsIC0uZ36nEhY+PtoycEd1JmsR2Cee555pDh9IiOZvzbhCb1pg
O/VdI5K9NVbm7Et4koeEXslTo9yKmv8YOp4886u9XAb9Fz+DNs4papbbF83RATzZiTSa+VCL+MmZ
RkD2AGkgLCRbcx2nMxXYyWSl3RMQ7xUWq6aJAASf/FGOrHHzch7t/8Vv4QJFtsh0XKczxo0W2okZ
AfnaQUL8GHkwf6ivjCbqLnBpBfUZrAKrCMoD+ZEY4WcdulPzfEcY6lLBdL8hV3AsyezedzXqXBth
g4KuehmmfXOlL7xOnkSAL+svlWznI1rq3WAPQL6RmY1kesbDYwATqLWW5PVYhWS0yX8WoE9xIjmz
ZtyzrU6AyAAU9Pd8MKRwgmuUaIFfo8mH3x3Dg7VPGYz8c4yNoWmzmMxO+qlHYDy942dEel6ubHbO
Q7DRpAgvQ2Jep7UZsdSoZtdxskRCH/de/LiJiZcI3YJ9w2YBAjruBm1227sZwiIK+yxLRskqw01j
HKkO1/hnyZmq1XV7WDtCnTRSOB1jA83Jx6Q12/Drq1vcNa2SvujcwqtK68R9JBtF1iEiRh8cwXZ1
aRWAUTlW1DkOcXLbvY5ruQcZ0n7E7be78+oRJnf6HSKqDSCigC8qWOKvXcX1EHP5BczrsDCFtx9j
iKtDT8iOsUnAhR7dlbaWhhpr9crD8QKyQJAX3S58VuxnIIZVLNeltqoGYoncbyKqZha7qDsdHM3V
Gui+gdgKY+oWM+RKSzQHszKcwonJ9tbT8ThZ26/ei2eGRd7GWBJicocATp+mu7qWl9XUPVhfWoKG
e1W1cwKCduMIhSF+MOcEfqhgaSJS8+2um/qvXRudADI2ogJWD3m69VnGjz+7Ak+Iml8qoVVgj1y4
dfHXLHyGZhNc7fxJQ75l5pGDwFRh2AYCeaY9lcotJtE/y7Vx5ie2hwnwjEic1Of98gyI9aHB0cSY
iKkDl3Bze0pCCG928YbShmsLaSBxk2RJ6nnuBR6KiEk6vlb09Ty0PDR9EmkP3ufsoNDUCSHHstnj
93mOX8d8V0c47O1EtJwaeucqoavltq/bamSv7qnoyjzmXkH4qM/bGvdHVliaNacAB996waX6K11l
TdUmYi3v05zPNwrk/bJahY4vyYjdt60hkqQNQaWfGeVMwoZAASEujZVYU+UydDI0QlvtZ9iUB7Gy
5q8scfA+RD/hUQkw0T075miGGn+h0RXBd13mGgYe9xjZdQqMYmgoiP/9qa5vidKUYVKuafwlXfqr
BBJ/vdow1QrpgUru7QT+Uxr/cLVN9f9gpjrJLRi30nRi2kC1vqV04P6F9qvnopqFKV4O/ZHVMMC3
eUgQQj47Kdq0rMDwqnRsvvuyyBCOTNlE3T6AADPo2RT114V4SY/gqsk1yX3LVbQwE7DbUBWhe5Y8
OiXmB8NJpHKwPNtmzh4/+85vjnEMsww7imGRH/FWdLu+hxaPS+SLFQzRCugpVrsZ8XKxNnBqNohR
u9Ecov7S7WzkHfoTQtOuz/+URVGOGOv9Rs768G3HC6EYMTl/sX+eTkEbJ1sZ2ylSoQuUYNLv8aId
WNywIUQGjgQBjr2Kqna8wXPE/heiW8l+wOUcxUfA/nf1RRSvRFvhy6KSMtwaiV+yqEwpuJOE94n8
AiJBanWY6dVlHFjIprfzVh1TTyqBu7GpmLyl8VZ7D/k7cnp+KWzkDzQfGEJWxme9W6a/hDpiyHsy
FZ+O+AKnJYCeAkGhCJW3ufZTAP/rVivCsJHIyZhwZhgPZQCi9fHNUnvylAZBB8DYugOukO1k7cjl
Du0waEiv0LelB9h7pa7qDPmDhJ3YuT5ftCzSoNxCpeGQo7c1Mufd5f2yH6Sp6lw5dZmmsmhSF6Ry
4duoaeX7ysazPLY2EqniG3UEJ/vvrwZLyfxG7ZB9kdVMELLFOCPtiMr75nZZv4y3nA9Sg6kjyPWE
/jd9+5hLFlBd4iCH2anVk8r8gNakgEfRwtDI8KmCRf8Zbpne/0fOkriIadL3YRX6fPGsNr3cLsV6
rJzzETRCvSj2yB/kWGEeTMTONrtDAHp9mg2ow0OpnNMH6me6SLHbsvU+aUDerqfw1PJt1yKoWPf0
9TtJggll5s6wdOjvK4IY8AsLE2T5130yKoe9NwF4OYPqv8qxgYVFgI7+BL9JPsPP1YVupIZoiW1r
jDOiMbAl3WCDU/oDdOswsOtyeGBJQjqbGtpDRlLydgKyrOiIfm2l0eReY/UnKQoxWuglCuHD//em
wM5zbRB5/qTQVU78cPORd1xwLkInW7SXmvXmzeSEu2ISC/9ZojeqDjK/HIbY4n71a4YF1ctwjTvL
GMWPcBipikjAZY4OMYS42ek5paQdttYCv1xUrb1owkn96moC7RrtlsHz/2lG6h9V+jty0GLlzNwl
8vGeD+DuMXfQbuV6xCJ0Yle/UqaPr9OBBwVOgGmx28vFDQ9zaCJPYuhT+eCowkQHCI7yNycn/3bg
fXHtJBuOZhe0XGK4PDGFCDOZbDPOzm2ui2ThvXlrqb7Ci/2Ha87IaK7ZT3g5pYVBA7xXbCCy345G
+qTvKGNYTPT3ce/dpwevFMPUKkECr/tcFFza1z0eaH79DiNcCBYLPY3P0VzyoJ8BVLOv/lpPt26u
s0UoioNt7XgdYGCNte6qdTQVVl0/qI2+xiz2sOXIqOhSlTOPhFju1rwMId6/2t/xhpaCxZsdGXmE
dgF1muxXQhDd895dX3+WU358l9I7VMCJ+ccVeniYVg97EyrntBXzReBLc6R4qauivb3ctOWR1E9g
15+DeHQufSYa0VDJlsXbJh1eufvZa9AfYmRsBQgcxWazsbJ1o1k+MwsgLEIGeiN10spPGjbMwree
9bCwox75BaXcx+O6B5LH8VAfnZwWWfQ3SxueppaTwUeAkRLuiTj9BglrvMuAsU7As7gWoy01hGTv
E5nfl/eHrZktZ+AWb0u+U9dOUOqaJlsF1+fo9BOEg8+jT+gY7C9qPLNApZKkijiKQhvcnQzdSQ74
AneDgkZ2BPTQWaHSE88tf7nfnSwrA62HEajyVJ7C+8uoPS5o1LXtn0bhdGPAWsadqu6iL9GWcwLe
1rbDTKnvHtzFx9Y+Fq5FJv9WnvJj2fAscyIMavbLAwQB7/LHQv+UCinxzk1Mdc46CtZC233x9F/k
BhgcyUTO5sQ3w9ZEj8WwyhXflFzQFTNSHnC6jbyB5xvcayxsCElBrgMPixF74IcawjPLTBZLSePB
mvqflU5lxwfrjvsRvDPjEKE+l+ryZXgpVriszXCkyBiRZKwl90lqsNkIt4tz8c9WNFcd7RuPyTjG
Rx8aT2Wbe0Cg58UL8JMWGwm0iWb19Mr+lDKX2f0v2+Pd2bxFbXhrObVii9l73gZ4muva3NXsWyYA
mvGJa25WA1xvHVYgDlCcNN1U/wdASYDKs3CN/34euqnwRGcKMGENkgqu2djE2/fuRBkOACe2A7e0
1vRSRXNST8mYHjw/Ihc98ByxWqYxuHfUC+rVqaejdPpiJWcfKdg9F6rw/+KEzr2G6KBKJSfrZef1
EyZqoALQLyJSmD/KOwX2eGgae5P1843rsVGTiu0AIElcG3Fgh9SKmXkYT4FTkK57C3jNpD71PvrL
5UJ1TgOZhlSXfQkRVuXHP7NM81RLnoQLcVraZEJC7cBLnctjmcdT+Hm6sDOYjv5TV5LxxTUf2xUs
StAFqHEvikRXeZFNg9RZ9t13yAm3cDKfTWaWaMJ4H76hkq2GufYan8MFqOynVFEaouMtHMmquOEM
PMVUaAeaWDLuafIvcvgVczki30oq9V9CrtM48+fYRw0BSJBiCr3TdauGyZxmY4oMbOt2uwAVgspJ
uROPhWMoNC8M40FWfpaTJSJqVAXuPraSHte4FrKuE8f8m7Z2PWgsSeJMGhup96FXo5BNNuC7blb9
i2SmGc9jcsT77jtJzT/zJ+A9eCN558R8UiKU/J5AIlcw651J6khLgyVINgPijthhKgX6dFDO+8h8
f8027Q2cOpLXYq3UBtazK1ka1cB4t2QK3EFmwg2X70/hsMCimvj/JzppDCvlDYOhWFOWLfErA9+z
jobCqurycpxn18upxSe7ikxwJKUUMBsnev150zWEJpSmU2dR5AJBl7rwQAw9904ca0lZee6lwrsR
b07a8dn7rEQk51lBa1qy9QH2sNybYGtDzU+fO2gdbnBKCHD3Kyea4Mj+8qTsyAtILEdw9gGebrjS
WV5GgcmP8OnKP9GZmupZSNq8mpHRcQNeyLRePILuU6RuQwUHDwBhugPDNxu7iud8kIb7KXSCUGWI
5h5Ru0Z5pPHMr/rO1rnBhdeGa/Wif+tdGuqmmNgBBLDdZA2HDOmk+vBJgdUdoqpLM6vH8k7FoDo6
nfEFkC7Z/c7Lg6FY13JNYG5xcTl/SIcq5XKtoPofhC3zjWfvWk0qWaBTkyoFLX3GYLXX+DcPHFbA
v66buzQBog6asVi094oXHa2bNOO3DtflUGOzUXZU2MPhlI2azoKQBI+KTXbL59N4d+BV4EFV4xLT
sRZpvViJYhspDW53EwYxctmWDoJb0YWUjlv2pFaMHMbeYSMFyLSpq6jMXOasgaU+QUsDKsMKaSnR
H8n/5V8E4Hyf4imfXXIIwJcX4jIVmaa8kSep3aI+pxqS2/SE9JiwIs7MTEdoFzQ0C5W6kxkhAl9p
fy0hDyC4q3COPW6I1oq+BDvvzyhOcz8fEYHaI7Ao5XIWN5HNWVQ++epib01sUZanjLzS2M81BMQV
S6MkAEbza53FiOuMZIJ7a3kG+FDzsGw9eYSrEpPE06jlLwr+uC+zdh+Qqk2WDbQ7TKM79Dh+90gA
a+MI9uLOlnxdhDDf74/HDqx8lqY/YdJWSmSpScvzXSrf0JQSe8cvfaCieMVa/BUXM+1/AwjnydWx
ximaHxBKMg7rdoaBld2bmLoyf4kiCnhrCBgPQ22ove8zBP8q8FEkdQt4llBe2Mz3GnJcBq3wBzL/
6vqSkFILPeRkw3iYoPfTRsI8kgndgWxMMkCYrZHLK50P961iZNY9zKaEpoeNnrjKqHIzKiGS9Jsd
q53lJKoG2GucjT/96SPAcWOlxYGEq21QoXzffhkF2AIupqZzLBZyVhqrIRlnz7wlxJhGzD/lLcco
yhq4qv8TXeXHXJ9ms1ZhbJYkZuX7pinyagys6PgIb71+2qNIydaeDoSny4wWGpz94NIyh1yvi1R2
RD4NfekRDalNWyzRIwFpTq7pM2HEUsMC2P8RkJCX1HyDFHcSuy10PKk5uWj9nlWoSRWNQxN3b7Aa
8irLBllohPVefF+5xkG3H22nRFduNY37PnqzTsaOSdQ1gutXTzGBR1rkXoqWqSV9oV9d8A1vzHWv
9HCpHcG+SxeikwURtwklDqDLncRzmfU5/YK4xCbIEAv7RcbOQAH8RPjmGbLX8qjDKy1DTDfH2ika
QTZM93FWAf64ARaiONRI8TQmwX98BTV3jxPSX8xvhJWURIOETCQ8DuqvvH0hE3FO++/eBj6qAPe3
ebGVbeNpbFQEymXfTBwJ+7JH6tp7tA8Vyeh8unucvrC9Q1B8tNlog5x1sc/7kgbOnSvrZc47ThIS
tfxgQ0Illm3Hqcl0eOyPaLTK7U5AycBLYk/67jDZju8M9jQpVoA5Sn2jhAtLs79H4p2rNF7oECMB
ypVndLHw8OzqSh90/nXxmsuxfQGhcWHDTP9DpbwqiwmbWDTtKthmrnIfLe3mw6qzLTVE2qVJzNoI
JWcQ8nfw+Opb2ZpmTC4V72DN99VgeG73c1g99empl+p0LISOrs6/X8TrdhxezB+ly0gZxghKwzCD
rkBG3+Ekn5vEY5fULY38+zMbAuXmj5AMpa/69VIIq7QJvpuNqB0o/N3MfG0xapd3n3vHd6+flLIE
vqkT78fx6Qp6qDnMke1hIUQWoD85g3wZg77GLJwtYCadSoLOnu51FWvbMVBvlgkcMe1GL7xWL48P
HwaAs50HrE9UPXyPOVIWExNt7nWYxSR9txhY2VuuviiNvVhh1e10xtLQGEpF78BO5nopS9JqHfzy
QJaY/4qiJ/Pc8vwXZBiKX57BJExMaFJ4b5FlMZGxHVXjYqCM1ffWdCwC4LFSiZQKriui9y8FRBP2
wf+6OdahZScYK/NCikEQjsZKhVC8nq1ATublZsc7Zzh/A9mm/4XnJqhmUyG3hznV5ukW+Kmzvdsw
8KyT3h3z3IG/HRnEqgp+5ROJBcY3+b3A6XXG4auwaTvP1fGvZ39donhfSxwSAoVkS6SFYc3wMfQY
Ix+szhueKhkTl+EMm2EfHstlKRGn90zSgylmgfYuF1QeZz6SV/amsdKsojfM0NsVsJVl8RAiYj5e
Ek8Wfyh70PSWZ8OaMxrmpPIlx23+7z5eM+e+tvmjQUPizy9PF9KxLC+YkQEiVH9DxQmIlDTiJerR
lv2hJHPkSluh3Cymv1+hMxLxUtt/UU3eqcTXkWbwiMdVTL4tXzW8LFhbSfjgCPfc6vUsAxdRvRbT
YxbYAGQWVLJ1ATDpnw7arh+foqtHkFo9rVGjmfLpERQDgZ4v+IrvAdYiC/y/tCJHp5nv2rVPJz/t
BnDT6X0yoh7JEw73fPFZ4YcNNwGQPPELfSH6hlomxDkJ37lTdWrhQnKTqPyStmK823aku25zlJuH
HQNBDAYDLcASBbsMw6zEQBXN5dwK2ICFKospkysZvCuSB1gdmYDU3sO1izQkVMazeiz5Mjm2ssIJ
H1K4/bYi/W03QQLpQOxOb2F+XHv7kH0XP5vpbeFIZmFttAwKLsPswbl3YFZOHdA8G/iu+KmiYk8Y
tqEf/f19QqoU10ElbvPEDWREDcMME3XRBd0IzcEHL6Ko1mD1pbSHFHveeXKL9IrtYhU8mfFQwJ8s
veVVGIxmuBcSKKwxPBjRRHd3hc0iODFBKGVEE0kl7QfLf7HXf2ZfusJBUAcFoYFdWkeydlrAu+wc
IxpJfXbmCH2NML+g/ijtm6uhq/j7F6kAKkHI4mAO6ramtmxowwceZnZnJfTd/vSBPQKklfHjJfIa
WUIwvaUz8EqTbVSrR/kFlABX3GaZiQnhObqI3+I+F8n3DU6sJLRvi1aWc9dILezxlV1XoO4B/L67
L4tc1su/L3aAazZ00ia2p4fq425NYuhLfHtmAt3feiHBbZqRO0fiv9XS/Al9y+kk5w/meTOEhdfK
RIcO0/5tCqwfY1ZFww4w0blvwpTR7eN4Pe/0uHU0Ii1HTOwM4sRvKq34gpcrrgktU7XA/EibYwKA
5f6hllzZA0r7L1Tq5FqID2GPP4K5UVYxaE5b4cxjIUFuEakXFWWQE9D/mxwiGet/HQ38yL4sQ/rc
i0o7YKAdF2VL9KT1pjPTBrlczlPr4SNHHFHSFgbPKVTTrnK5qOPJX8DzIUnVlfu9aYAn4BMNRDGb
m9XyKLE81m+TuY7T4CwdcV4oCMnh+mYpnIhQWZ5vOEaZT61voRYJP4C7Rouxrc5UhnHam7WgHN7t
BmQ/4ygXYiVaA6HF78waza1QdXnyAYt8GzMJ4/vkLnCZLKixMKXy9AbpXH/ljQZur9W728IRFVkj
iYLSr1I7/phpFVVOq7TiBN4/46pAPtGWiDm+dNsbeQLQwm4x02ID9OVAbIdjYCG7EmdmBXBKBSQ8
6BNHC/r9BzxJNur+26FoKNG/uWJwApHkVKzmJgfviCC4o6lDC/9PsQo3oAK0HshZYpid69qUvMWH
td2yfF9RNyYvuvoYjeT0dSkVQmcUo5BV2uv/xTcqz7nWrUlGBGyZOxvVZ49ZOpPqtlHO5dtJHp5b
+Wr7653UBD6Ui8ExAgL170nUjehawvb0C3+GrmockeMHYL15vElyP3Po7PrheDmLVJYFr6Vn7clM
PvbAhETi8JBEq1vvEoUtVBoCyu8WN4WNfcT658hqcNBomI8pGMcSmHphSWWieDTFASBECXrqxTZa
0LXX8Pqj0oBfXzbl85S7uC2DxngIf14Q0fQJUGS4xF0j8klh8yQbmpd6/WKOJJLc2cbz/1DM6Iyx
+Q9Y9/7TCGxQAxpfFoX+hWuw/uBWutejaSNbHE7ILaIgdUPGuTHjh/+5HGdO6Obg3Is2mOvufg8f
Cg85bCb+Llb/xtEtqfyANeZjBs9ATQW0maX7jsQ+SzNv94axDjaW4OniF/wcV16AaNDWXnvhIBA3
TCoyF+ltLQiV/lT02DvOVetAwGcJaRStBQ0R2r8Fce5nH/bAKgPHRRF5lG+aDQ+i8mqR5ZJOuhxx
6Zk5B/AD4OzUOlCbBFzeV3y/4YIhGYr3Ac7S9It6zlnHg5HYt9ZSeIJvbeLdX/niiaBSn05BPktv
F/fCSxiu6lNCmOu5MrlbUZbE8FqqGoSohrai29xVoTq9S9kZjIxp8EGsQAXZcCAUtIlFdNiORx50
29Fig9IB/lLE5OgHOjVmvmEQD3wjQu376mBLlDWgBkO4JxlCuWokA1em0XO1mdoVR8P4uqZU39wg
PU7C5j6+Gznk+Be2rflIOFdgSVcb1aQa3fQxME+jMpe0PdBN4u7vq+2gItrQ5JTttPT6YdYorN0R
pT3PSJ70Z6YZSF2tBSl1h2hIEpyvDIA6PmgBNEOrBa0Nv1rtvBSIyKbsYT2sIDqQMuZgOy7bA3qa
BS2fRY7wLLTA3XuKJj3lkCmqq+ebY+7RQ04kXrjElDewRPSuAKKniMpUVv1kLLAnewmC+p4btaqr
LTQKeoJkYyFnUFLNZdI9CVlXs5y/oDSmz7GToFMEfHSOFGDpjftfaWj7JdVSHdNWQEFaE/QMAm5L
uI6veg3kU0Ri9CORsZjjrBIkAlK/lqiCH1F5zXv+rpaQ/4d/F6QlmPSncpPiGeJgzhLRGzELBXNH
sX7SzAh1qn9c07OvE8+pflwAVf9gZn/gVgqA8kv6i7Jv379HlguA0/4viAtQuopSr5+HqgYl/a4q
9HhUi5MBTZFYkTzFfJrEjarZHQpoawkLvr0t9u7Net0CPerTNl2Iwq39zF2CEa4oPfSbpaShIOe1
X7m0NBwUOnzVisQQh6wTaT464FOL4r9e6Kn9/lxzW8QcXxeArp6/ORJZ1mKBg09CG/bqJny2PDlT
H5l573to0vOpX4KFYNx5JVkLMSEnWbv9VCPY9mLZYmUM2TBO0IcW3cIbM9xDOT03JKLmVNF255gU
RQNy604HQbsSIJD5sQVJoHVzxy74ZatwS4aAY8eRMM10UatMutbDSdAqA97Jp6Tx8WDbAOMhkTVu
AJxuW5PXQHWjxW8zryyQ7JtI2dh8LmXRYWPLPfb04SfK5sQoWFMx3CdU0BdxZXWf390DybPdRoa6
fxE/QodtYjXVkHpEt11Gz8KT+CHKdNjvU2Kyp5/KMn0WE/bywwdl1HLWgSAzcbZaptsU1MZB24kC
CCOFL3vhJzou7WjbRY2te9BA4veGorY0DrVOq9wZjJsxL/P+vvE7AnzyOp/MykM+yj3Rvk/tsQxg
OrCQ2EsvS8or+7ZguDot5N8sKG3+vPHlXGid3tCAkb28+YM1UwtLiBP/AkWjEr3GwbnoKokmIQJZ
Fz+3aPUptWW9E3nrY2f0tBi/KN8bMob+dAoO/tOaeM20HGGx3CmkBUJR1E1GqrYio88Wgvb4k/P+
IaAuGJvS5zXJLXXBKEtkYVsanbCJ8mjv7Jb2ah7WB8lYm7ctKDRydpZuTKAqBS7iMqvz2XgpW0mG
8LjtWVv4zg2wMwUDPS1EqJytTAEKWVvhcp0dC+yd5oWdRkW4G4DhJ4uWX1oahFGnfleykRGtYlxN
4eRQyudsFlN/UQ0gkmu+3Jb1VhfHDDCiR5IFQ9x7D8jbtuXHm4hvHsHvvW1SMKSy0HSv8IRQVv/R
B8xWd75WE4llfg2sSwJJTzI7MpcsNS5p2VTfTsZ1tkNSFLzz1Lsmyjhu/76jAGK+vTL0bTzB8yUI
gAXrvhe148echsNUO0HuARgKfHdW6Z2rXr/DT9rf4XP8xzBpNkzItrajW5Mv1z9/Bk5RWLKRl5rr
aNS3Ytwoad+D4sgu9kj721d2wBd+5l3ObjRE8si2s//1xjP92XYjCV0bTZEWXYjaGKes1knq/byz
omI2d5hoHPxdrJ4K4jwCXw6gFT3Z32mHpe4SYfjtbaCa0+LJfAtFC0CD2d8uWcFfrOXGHKUrBSF1
xBS5Rzg+qUkH3Z9ZtVGyXcXecoIbaEmc3LsjdbRoarwG2LJ1FwTOnj47zzlDr8mXNfGuz+03+l1S
/Fy2lW2fuy8BOKKIhKO02fjgR3YTRT3coc5Xq++n7ID8ehUzy4L0uUyQPfui2XplSG0Mz3+FOmQi
yp1UE5ik0g0OtLAsvLCGgVTDA14nP9eAPpnjAScy3LRXqCrN3/ni2GdnR4+pCloAv6UsNIZu9o9g
M5p5DBGNbpNNkTfjNgJAhyiJ7zYqO0ZU6HG/61kqQ5z7PxaiiwNnJBEF686QL907BZdWJw66D9+c
cBHFdccem4acudeD2MJxE1Zg1oMwi5eOQ3GRY8903B4PhpIQWPVlS0kgSsSWQnfcLeSLM34rzW4N
jkF6tn/5647saRT0SRjY7d1s25rTw35NAfsFX8cKj6MkOViDu8sveVFlBPtV0wK9KoDYM80IaAoG
2Va3CA5jy3J9A6XoZoVghupokipsNBHq2kL6QQPNwwkoIZ8Q9Z12DZR1V8uMJc5Ri/LiVj2SEwHj
buez+dGiAvLWziK+JfPd816bdByUynL0sSYwYayFCOQVkFyJ16ogHO5q1VethXMQqfJVtD1Iz9jm
nBk3Dl+8FsAWOIomT31qC+5qMcosLNYPfkXg5XjdSGIoeq51LE2J5W6GE4YzI2pw+P2B/mLyKb3W
VkW6EGIMQdHCo6LZHI4NQFXCtZxu/NNiKg9UoO/8oq8aLmcW78EyTD0q1ly9w35Z0M/+r44sgNsX
6XmKqa0oNeOYBzqHFM5upLrzvAfuiWQCtd6+bAzio9UvCnbBtIpBX4hpeVZOp+TCMjPQHt3p/ffe
ni4J5la/hLoJTfd/UsA0DyLfmDeH+5CZowoG4rczf9Ec7MhVgfc/eN15hEJKsCfKOSv4mGzQFDLR
GB2t/AlfnuNlP06asEV8SwAA5++Xl9FxeleNTHngDXSmw7m8u+xHkdRzuiqyvL0K6bwhLvb9dwJv
lur893nLZCznwcYqnrIrakqkA1j2Q3Sg4tbkvgV1ndCSlq3e9V1dmlnvEVYgxsS76u6esoJITB3s
ylQL4LSNp1MSYdRrpTw8eSP9nfVczAbqcnXX24cFA0efX7ulP9+kQaeWx13OOj9m662CUgBNWkph
tXvG2dNIIvj6flqp75iGM+SVBzkmVhZYOoOZhbZnmD4IN3TDi044FOR2TWLT2YWmzLFw3OBTqTCg
4LkY2FRF5zSXBgKQaW/BwmFdMMpWHVTM6AVMu6J2AaUVBC86t0lp5sjunAj4QkB26f2zQc91cmwY
IrNF3gHju3gC3pHtCGN64ml1U9WL0G48O507x7PcfEJxCR/P01D8Z6+Da/qooRy49bjSS6zoefJa
+WvqdMYHFKUPJEMa5MWUjMbC8kgyiBfX+PABNPayFSQ9krozI4oId0JQlzqX5gbXx8bdbPyMmd1F
fX1v2ti+8W6z1gSSO7SsHni8GvIzetUlJD/+4VoJm8BwZvn9iUMXX/jLxG5WExL5E4XOX7VB6dlt
EFHWSy2h8YoFt5OvnQD7kNEfUY3UxrRa1VxQi1Dm60zdUd7wYJCbBj94Cc+oVRAHLbJYBxlK2ZyO
MF09jRlh4MdpzYm9WXWT6zdkTMMIxpWqyqf22fA/QoXl0w0K+H7vqmjuJmq4D57GFnS4ibT6REHK
1yhSy6WbzkBXtW71GFGFQ8YuD3zOtSm1vumgqT1b1xExSNQICmXHhftTjj85frQfy2FYXz2mWcFQ
gNb7OZbkenO2mj79iGSUyl6Fo9L5yFYpSDbp1aXpEKC+h2Z9Ua3ParLdus/8LacRB1La5CQiskiR
9DQlDH3aHhyr+pxxyJukmNncRPozDS8HOIbJUDq8Y5GfyOAupvrOeFW71925dGcTtZzEK43qcX+O
nZaWc5XHpG+iAmpAICRA+AIa4gzwn+WIsYMAIqCVcoWFshq1913daqhCyinbG2in5Hybk+2AwKqG
BS+f6T8Z7Gi67InILTR9An1SW3ln+9OduWQFkVF7J95CZDuAVV0KQPcoZKv08bJ/G5IAky3cJIOm
a1uU3lxvIvYOaJwml0TMCZbjfNuycYplyrFOMEpKuRDRXExbw7dA3FWAtePFDkmhal8qHn74Wn2W
VJ2WXlsomxb6/wREoLA+mYkp+7VtQM5nON7mlU5vI/28SOxqAk3Um9Jk4Q+wcXJha1p09KiYL9I9
+QzYSxXwxRqFRzqUki9v06e9Pq/rISuDSj21ckU4L9XJo3A+8uGI8fObNJtxF/nkLaiTD3Wk4t2r
YgoXOqXJgwRc9WbzA8dW+lg3l4//Zntf/UkzWSz8orS8dmjiC/COeso1lZ6Li/KQdtnpFpnUya1D
3KDkSWpotjXE6cXV88DLsrNXhxGiqHR0XR2rSQkJ3rIxehXefUBKB9qHq2qZ/deSDCbdBBxuDA9j
hyk53uyCgwdwOHNTM0xYuORek1zzzu5Zr0W1e9acyitvimCEmJFMzFdG0RTuf2/D7wJXKgo1xL8D
OEgj9oEdLFkIE0A1Ypgrm4JkYaGtFqRUXZazVr0L6u3BCqTRVDYXLxZ4bX85WNQ3oDI0wafdaDnf
EmLWkea9tBp23GK639TkxFWai0BCN+xcgDC0BLCMln8f2Nb9mDyoV+jyg/Qpg34bQZOD772X9nuW
EJI7s0+hCrAFpM5YtSjUF0zgHyIxh+EeAHrMuXkXIOXhdy9vMhpHAkgqBDO19o2WSNWGoZg3gmz7
QSDga3lpjoiCBcBvCbaj5c9yycRpB89ljhMMZDxqCrg8zg7R+yy2WuP2ee0tsjZETswXaHaU60dy
FCp9yneX0di/EkW01oQ5mqaZN+pu5WFUopfc/BhhAMQteJwemvNCK6IJ1acW2jw75bOr9us/DZjr
cU/zefYmWCH4pyzm31kKaZAjdLVyqAuMffIGF5qRmi4qeTFDp9mJLfVibQlAfex5xTlq0gDsup6o
8fsftRlDrmO50xcn3QDpTPWJNcC+xZN4aNUyvMBMcUOZdUDHzJ6f+aN7CeZlgix9F2GiN9gH/PiS
MubrKCpxOcnw/fjyRANwgKpVs+TDvGoETGVUfNRr/QoNZ7wPLSgIN8kxJdZ2tJF/CX0cnWlRKgQO
9qzoEdoBQMBAgh0gLCSsuKa8cLSOd4GCEYmmYc+LvLCJn+BmrppR2NY+cQ13vaGsCDAxqQruwbky
dJMe0PnnU9PyyjsZR0p3VH1x7urle4JiZaNIYTrj+r6UKn+3W/ss9jUr7sxem0gbHc6sl6oRl3J0
MkyjyIQV5l5gxu/Y1s8yl2zK2iZRZh4eRwFWWEFKPkxMD9OAB5/Gg7qunBHpl5L9B7UfG1ub2lpW
XuKJmc2fP3YtXZf5ygHydv9UdPDrZuq0xuzWhAE2PrajT7XOHRPmklsw4s9OdmXhE7WeOq9txiBM
JU2QzIyt4jmxV7HzoCIcFJgtDHCPsBWbnBcelX4/Y9MmxpT+6XlFzJvrCrFsDdVHiuY9prc9dOkr
ODiPbz23eZ6FyselSBCckAcumPxmogO/TCR0YtXTStnzbPS5Mls8ekldO/3BeJuJx6S/OOXt6AmJ
ty7HnI9ylcJy4xde65hF9W9DEEDCtdKOEiST0xwnl8Mw5lhxMkKQbImSt4sv6ouPHXxUiqFA1iMz
nxiTYi86c2LoEnjBjT5a2wRWR2l2uemZKi+QG33w7JX/2d9WMuVUqCMW+Lh2WGITIJ0O2F8KpIU8
TXHZEDbQU9t1FNSOs0hUI2K2Hi1rZWf3KO+KFXjAA0AdOL7UVqA0Km7sRvG4oUr1vPugEB0Y13vQ
AWfjVV+IZ4GuU/etKaM/WUhH+/PcO/mWhtMjCVtPytE6vX4MAbIQleG7eAFEVfwer5PDX7PU9S0X
vznJkBgp0sE5RcHQhHZZO4/e//NlTfPB+KNpxA+rwkOz+Pzbm3YNGi8jA6gmK1Wzd1qgnitLF3Eb
KmRwmMz1NU0bSDrtq40Ld12/dC901ezpkxJnEtxOyC6cdHYlbTdXBEpJJerkeMnRcjVCOFfRdeLQ
+uWADOIgL2Z72GJo6L3GvcGbEtMsaOYWkXjEHhgzNxv3hdRhZA3L3sJwBzX9CzMbgJAtZyHCCfHM
rxXecbVCgpcOmVsNFIv/D69ZlkOs53LeaqOdk+SWJE40u3IqqU7sY/jF/ifglba9pwtTf3uJuMYT
faPrcNG/tMLBFbX2ntXR2LMrGK4Q6Qwxh8TGcBsbfKyfhJ/HYkYOZ5MAR4JLV4XzO2xxhlwoCKrZ
tUr12PuYS26CGVcb6ub86xaieilUSWwOBzupWLnaDAsxOkWoJWS+FvIXa9NSCHxViK7ZumxGhLfs
rL/UEpAzDljSWawgdgxhSwjaerYhNHzcn/JcqORsYlglfYEyaGZxWipFXUque2x20+6GPYQRCDIc
Bv1K3eF1PpTApxY6SZZ6x3/+QULX6eEnxb/pevKvYvj/5R+9142SCxXdgGE9EM3NeE2Ty0evMCiI
M+9oEQSmrk8K5bz4YN7y9bvS6xw54joBpYcEIseb+ZJ8plkLAWoMrnkH4YRw9VccT+DInv9cqBeI
NYh4aAKsSF5v7IPN5t2VW+ZQriRi/hR3oHDeu5JIUs6sPVALnIc0uZ5rAo2Ti/olp3OVasb/3CR8
g74Hgp3Pg0TYfNI+Yn2aIo9975Ucft60PEmIuf0NXXYxhKKNDhDsc35GBIqdxVTB4bsgtYhDdS62
Sup/YqmW8YT2yCBw8VrSfhxoIDVkRqD9LmoxlecQ8Yp0vgQS4z4KmKgz1XBh4v7kO3mmZRPH/6eH
Y8pH6GARLNkwQh6FXOGeY/Zt1qe9HU0GyK0PiwMOq0+IS/TCUIQf+hRiwseSdCa2I6wQ71wGgNXZ
EX/N0PFCurjlnzfXyXXOAoSVzbQfEkcvAmKy2IiG4Fsh6Ae1c+EnirBo9um7Ycm1aqxVDzvWLKMm
iK1LVYWl5D+Bg5WyNuu+Cg7zmhkEsDeTN+MetD/tc/4359me6z3JoKCtVCR9uiGZafOUyPlNcsjH
y+8Z08pUsI/UEefD74ed+oVyTJXxWT+UEpUQp5/Oq3aQ0FvvKiLum5F7lnzoVBn4vA7zzPBUZeeF
hLzLOyG5jSiw0sautpLEpw8jsAbocXcgEvRvAnQjiwXeRt9etrc5/9lVMDmb9Ks+XBQbdbxRxw+Y
moHQva4wsc0fm7ZDC/CulZ6+8tMqvIpT/a04RRyTC7b5t4/y9z4LDhf+m1AccwAiq5f2VxdgD85k
X4eSMOrpOw3tPzh6KSsKL34GFhVWi57SPMzv87e8B2VQisDllzEeI6wTD4Ycc60tcrmF/ujO4tml
sFoosa0MMeL8ffc7l0v1uS6Tm9KtLQveEi+VW86mGS0Dav9+bhXsvpTdIPa6yef6aCmY5x64FgES
nwpFB3CCi7VLUckHGyaUiLg1hEi+pfUWRDTH5c4yuMuevFMrDGFRohsATAg1rbgHR0Z+so0LNIVl
c+IUy63szkLBHG1EU2RHKc2iHEHEAKQ4qznXxS9xGvWjvUnf3lozsH4v/OhtFEWIulmpMksS7D7H
JoDdmcJnuBRyHgbPhyXJ10Jjc+xR3lw+4k+pCOlrs6fqKycdblOP3K/2PEcJ9r5ad9p0x0IraUHJ
7tQYRRIQT2XWrKduZvdiBzfGcVWgy3Z6qrhwpzXqkqrcUSNIYjXUQ6Vohjs6hQQTRxADav1fr8zu
La2GVtXhB33hPonPZbArAIYrjbxEl+Ce8t8ogrzT81+O8HywvjKF9WZwDfKhHdT7q/Mzsnfwmwnh
AAX7XPhuWVSLf/kSvTA4nrlAFFuMQMeQsXR3qt6EXnb6tuWUeeZkbbhP4pdVYuwG4ASydp63HbCx
C8Qb/baRz8G4f4yVtie35/UlAwCPIi7DKyVRsauuTMBya3b1Q/RXexJmDW2ee1V5d6CstXRYAMpc
mXpcjBdu89inKp73Oe0lq5HfyyajwbawcS5oN9X4+1NGddPGP/p1Nqw1useHeWpYcXDuQP4YCKNg
s14VzC8TTapHgQ576PpwnAPj5uhi1oKfoxNdiK9RdNdzHyDolcAB33U01ZplpvoYWBKlZ6P+Ii2n
kGYnAqvOgaXCv1L/vW7n/30a0TKx5fqKh5lU72s1X6Rhs3/izWSAAuZ2iUFd7GD0CzfX0MQPfsE2
4c1BxelY/wDO9sfkqcKEgg7vM5VGAMJeyaF+zrXU+1fZlWJjthHaA7H9hFGYmllGZR0rhZD++xOq
QBpLbvYj63xKMPDQUY5Z/IgIrCbQz//aBSTimq/O3Dh2yNgIMykPcBT2Q69r0S0gulot8IsJIwPk
KKueicentSxQkCHTpeS9WIFnZEa5sPpqI6QbcQm6dFA0xqWxxI+vyDlkj5jMgC8JVYT+fMtpV8Le
25/R41IRsHx2ZBjkcbhBxM3ukYKRhdV40dqLTAc3cfXYDms5yzKGzpQfG+Ixa1BFSZkAZEWZFQ+q
d7RhSzMffMpFMEIIvytHbp0a8RIt0c+SFRjUrAu2dS7FpvLqrBQxAV6pXZfBS4kdtBKSGjIXAYAK
SIqM+G3E7QEUF5yMq7mn4OKcI8SKCC23iyBIpTLH1Nc8Thxe8EJWo5FrbHKynOC4sSNPTS4hDBAI
ZnerE6q0BSO5oIsNUCLSdfagreTDsCZcnQihgsEMJsGzu9DyvY7e8hfZryEDJuRAhXot45dkr7oL
w1p94SWQfC158QeSrxaonJgSL5TChnvYfOMijIpOMvFWZ0Xgc73chxVnzGQH6g/q1FGnLiVP7xs7
yELC7NjW5yB01BElFXpHqyzYTOmMQHc7ry5WBizhMJS0n5vIR5fwWCy6YW+kugj9XsG6IloGetKE
UPtR7bxMz8zqVL1zfroffsMbCJjSP91M5++82B2GSqI705eBsQbGbQMOIaYVR9I9R5V5CJMWvIn2
zvE55l2ULegVj7eugV7dZrxx8HjjsPHmu+0QcA7UF8WAsT0ZB5ZdEfgPUwcOx977Kbq/MSAJmiic
Z64ZORdjG4OZWOdsQF3xui6pgYqOyO2ES6fUocc9w/s1EaWPR7pu36WXv/hHV7L8PrjPvH0bM9rz
Fx4dklwy63+fkyOZjYSuVgiIHEOaYFAFVKuTUgsdDzcEjfdQF8zxKV3sBfYyLsDVHBK36uqY6+to
XKKnHwd5z+tEzajBAlzkurI7lRKjiXnF1YiAhnwa1ZDd0J8ST9N27edKov6a2mvpbRHaOwC+bw3q
Ze10ifvk+Ha4McsmVVIWCB1/eNYcXky1vMzbw/T9OHIHhXV0PXPSJHPZhKl8LDiK0bwgx55rRk7+
XkdECO11i8u9USSS4SHuQUckqQwUcKXxfTdiRqZoOWdHO9zHUKV+pIwLZ5h7cs78Ld/FxNxwtSRH
q4Mkk99/XS58UgQVLpzQCeGxyP/BNSI6ZMRlktH7mlj1YEiZlardUHWQOJcvv5eQjj3Jeg2VDRL8
Z/e/pEnx8uZyBPVacXIL5tGsvkvcbtLZ47ZV32bV78NXiaJ0KlFcYmp+W0a0pert6mkU2VhI0KWD
NH7OAvfuWG/xtj6s3WMCyhkw8Tt1+AESDAur+GdSF9MDrPaN+Bc4Z7Z9cXdB7fZwlpc5bPCgQSWp
2Q/JTysBcw8BVKZ4a377Vmoc2cJ3SAIq7qIdE5pOWmPUukg4eQne/oTxVs5306UmCSwIsDaOsHQ3
Sxg7jB3U12YA6vldS53xJxVtbUlgKro3ZenpjQQPeo3O5lvOsQhqtAxHseVFJFlQQyeWyLvM993E
lss0z64FxzqkarbG2OKZkxJ88ZiZSGkFSAD49MbqHdcrM24rDutYx3Zybcdp8kxtAO30Bp/leU8+
0oJ6Ui8URGLYsWrZQHm/by5D6q15xiITzAqnY+gagaZtGv63sBkxSUsL1jbU5WA3JvIUiYbuEsp/
uDAtyFhtM7w97hST0JnN3kD0nEdcGPgN+Go08fRCBmyVoeKkDgHYWEJV3T7R4uncJ2HZm/HtEBz1
P57FrYq/qH0HU0J/iWrudOGL2jl7rzTDgNrGOP9y1BiCDKMN1COtBPxKSPaaewdaOxO7GB6ybyU6
JUbFB5JrZFaWVxsUMpNufY2apYFy1LTktOOgFMFfeNAIOi2nFPh7JfRhzxAe7EW5OYado7A25M6J
HKLJYpniuLYHRmvTvGqAbCbolDemiLq9yN2YDBzGxDJzD8uwJkJTaHW3+Ns3aFanrWA6EmUlw5Gb
xk1NqAsnYvnaIF0wjMXbVDeCBlWcdozPwMelywvwy5caOeNEBK6cRJjGcJ0Ul2WK9XoxlSdthzh2
9wSOjKPard5PBER7QGjkYlq87q8dbPYPJztjEv8SID9EHyPkLthH+AoUzGQb8FGh11hWe88yfZtD
TTK56C7dclaZ5J9NbSQ1JTkypezTusuKjcjBVlCQzFA7mWIJS8GWWEDAnNh8ltHkA5kyH+VnhDc4
Q/vHNECijmNug6yx4rtINX4/BKbBTLU6VmN8iAnMat8COMp82nLgtH0pL5QNMjLstLeV0C6qqcLv
JkLqLRWrT8mZLooqaumcCPsHnQg5azhbPBef5A2A1Osj0pqzMMGNCiOuhyQQk7ejlyjYYx7A2jpc
STbSL6B+tjiTuj9408OyBUBWJ3+bJLb68chOPsySbPQ+giRp2VjQ1Hge7C+eRtqwuqOIwBTTCmqj
4Sf/lAOTzPhwW4Kuy9vYOjE6uPHjNKCtTW42ANz8rT6jfmax6a6ijZZiL7GDqmpNPrt4o27ZCrQ1
CPmgnvl5vj4po57gSZRbdVdBnV6vBE+lofiaqi94Pm3yMhGIlZ+Da2mtGkZTEn3RdeyTUYRhrc7I
Sdp7IL4P5DMnauxmQgCt7xo0ZTlPT+xcrl3eLhLcrdYhFmLWPaPmZPr5TEK/WS2p2m3yCEKALCt2
XZOwplecfziIuDtyzpBEvuSGIiBrS8+lWGVqVmFm7Ki30r4xIr8bVWQbOufoHNNdJSBQUUz7pyjc
YVyLjWhag1e+//MG57ewx+tsMNr9PcURPp2uRNVd+q4cp3jnhKKOODDhOJ2btIx363EAzWjWcS3G
ck6mwaLZiBkD+I8inHMx4WhWLCa9DEYhycFwJwrU9xoDLYTSn3o85CB9W3pBd+KIiSyDbfKs093i
s4wXj36gnZrwSJfI6l5UgVgHAvFRY1uHTwhmWqUMGVZL+vB0MXE5MExmV58Fzr+lEYJpoZG2syE0
9s2Xw5i0sCWHAPVYgPtEdKeGF45RASw67XLdUJggLmQt7PQBiMoXMx2kmt0gia6ciwowNF2nxCgM
/XrTIp6Ek4VdYR7Qf6pEbSLnWNBEj5JlxWxy2d8fZyUdGeTtukGXEsgnEtr/f19hvxj1ZpuE2Is0
o5+QqOxpjmDehyCxnib2GLZBpqBqKOt6aIm4x14KSdwyeAA46GPX59d97J6xy551cXr+3TbndLy3
RaQrqdMR8dxq9oMqr0WBhok936z5Z9+4xi6+ruS/9BLnS7DdDWYR1sU6unUtLgvlJehODoAVqZr5
z9YSFyQH14RuGUcrfAguq29f1iGO2O9GsPl8OTwTVr/2U5JNAa0FBMNLhkHWxHQ+HmVc4TO5uEab
+tbqaqiKL4wF6Hh/ZzBxXGXFs1aSDeuPXFo129DeUirA6vDCFssHuzPMcV4J0QKk3YL6x82gwqLs
MU2Aej0qNSREF5TKZ/cKipJmJpoQeVEF1f1Isw5/Mkw+SS3kYlzM94oYg92fN44I5EMJWHk7U9PE
H7/1uEslUMbEQAwbk+hlViCswtk16xZAJpDErXS7ZXbamYX1lQo1Or4Ct1d8IEfOw87UVnD/6o9p
ATUGs7TIPZ3eKYVofektIV4htB37/bIBzqzPmDmN7jsn5wi9a1IsjcclrJzavPCHtE8oG/KCRm3e
ecU4w2OStsXyZfB3z9q3YKIdEG91tOp/63hlpk9WLWvrTNr1nrt10mY6MGJvJQ9fwr82yVkVaZyg
46GGp2XI0gwjCblFBK9S2jrci3Gge6R93nDxkA6mYR4/NJy/udKTxGNK348wZK+SzBfk1eD0ignA
GyrhSkyGxXzMUUlPeGt3eAtADE0ITwJ5HSrgKQ8jdi/Ezg5NgC1y/a55+0pi7xmszeWGz5FPDkPw
ems9VbzQy7+UVkyzwgQ03vd9TU7SzeJGwzAk89Z6EmnQDhwbHuUlb9SU6LMYK0c020r7wOKeBEAZ
XYBvytIlAFZC4gMVu+scdFN6jADqmQviDFMbWArZRQq9Yk0Stjjy+FNaYXbSnso8QAHPDiKQuxZZ
ILg6Ova8klYxkQtA1zZvNu3x/1wkeOk9qvYnrdbWM4P0o8Rmyh13KtVkgBzywy9ZKpoD885A1oHw
LUYPDAYcX75kYT5yRUs80fZ0gjmmsaN3Fel2kwFptjoh8GmvYHR/IY+oXz6OXLg4fykMLzJz57gr
O9opPXTH26a1+bMVMwSUNoR8GG8hpaaNT1CsFOD/baARzmahvDSckDQPkz7kl9ZmngWBx82yGDb8
HZ7AitBtyvbBXkmiDCbOz1XmX2TgNYWbDCIvHsBWxmHIvfCZbKJPXzwy3ZwZtP4QbVzws+obhJco
Zjc2SEiVLvHQy7ysiaSEet/3HmtOwZDVbevtuovRjXcS1F1d8XiMdVI7Jw52LO0SHj1zFRXcvHhB
4XLiPnYMD7NfHHqgd6t55PFbJa3HwLnHu0Bmr6rYqMEclpk+vDrOlneF2BL2lKT4c/JiMRnOWHLm
1SM2YyHkT+0aKIpXdYJU13ilcvfskPlyIUGTJGcxg1ez67z80dd01EYmTT2plwEiEktIvycAbeS9
d9un4xFECutYn0Pr9ICXz7aUsSvlQTPAektH2vTQ7NzWi0mPVWm02cZq7Z6CtxylXZjSRrzOpoEN
p2r6tc08saJiQNoZ3t944Ga5bFsi5gvSxXx5dQ5uOp8/boRVlfr0hXU4gicMKgWZCnx3yJXNP/JF
pYf5uK8RyneRK48EQipzXT6una6heSS+lda2SGK28fBWsm1OHf8keGxJQRE/DnrT4Lg4oZCoph2T
/KUTaA/obngPs6fq87/9kGk4ooJhLnnURaqVMmfh5/YZFzXd1GeTpDNgELF7jf0cidUNLnHSeMZz
hR74HHzeYIWH7Mmpj7bIC0OUcpoJrmYeGMsJJ2T09Ivxb4oT9zRSNXu9Kv/W4SOg+/qmxyWGCsHr
vbHujMcDbAtWIfkzrwcxgZRQylVGGeXVnlHzEM8ELQ9q+hiKPrfVTpULyrmC3xteexabVNs9smJ5
+2gQzxAUfplkV6k37zk+7A7mEFgnBRU7PapHllHaZShcUfRnV6OL5NTkvziQLJo3WzkE9ev2fHrG
tQ2lNCFQLI9fos36j1c+adRVOgWG4FANrmoyFsfJoG4u5nnDx+wzpoMNag21XSPGHR+uTnntWB9p
jw4ZOCrDB/F/jAUC5NPRVaMvJAuDJpHjkRB1VYT5SCS2W8Ks5vtJXb2Kz1HMu5Z8HHro3a8SnPEv
ygYEu8A/7p6bfgRl0pYiGSZqVtAHGXfYTrDNc/t7fFiMJNpFBITzCzB0pLfXGkr64sXjMt+fLTde
tWB8PWsnIVu4t8S64J95Y6pjrNKqGqY4pi3yz4YaU/M/+6Owm646+1jOM2l7aM/ja9tqrx5RmBKk
YZBjaeGJHNbzIOekX0SooxzUUPKVanWL/HwoIzAP7QJFtLRCs3tWROdCiajqUZ5XvvrSXVBLIi0H
seomWCXN0bR3qiwp9+i0bqfD2OtJVFCumJgahUaII1pcHO33KbGzzzyXbVNHHxATGObAAhk1CRRW
7PMgU/DlWUk42DSMb9CquRC/E389h1JwE6FZDLyXW9CU+4mchOaJd2G1sJ3Vdm+NJ8UCJ99C3acO
LpkXMBadAl58iNfuKyjn6C7EkbrutyiDqx9GeG5rda7iIllZAc6ngCWbjIuW3gjzemba90OsadnS
oLR47aE4fpD8roZkxdFZnRECX2FIr21HtMO+W6m9liIIYJqK41JoV/evbOFFIXaBUSrN57/R0pKG
emHqLPARF6Q2apyHlA0Bm0MoO0uDnUZ5o7ai+W4G+9m9o3wCsLzLFeoSZIOpIuzNUvzTkI055Ua2
PtZfp754Z1eZJIDSo/Q+kRBbVPIK0IUk0z0iqJRMs7hrp9LVn9CeVmRQyYZiSu+DEEhapcEwtsJu
jvyGrMLokQQgV2uYwRtms7M0XdJlorUeyOruh5xzDi9bPpFq9GRv8I9FINd0J6zmkB9kpSdWPx+k
8GqsIROIyZ6H+v1AmcAtVQAh9CYW79ifu89e8KFTOhpfPYGioIqxsftaWxLg1HrDeaKyCTiwbdea
qsEu0xoGg987yPltEcA+h/04S4PPNZtdOTEdiUV696Zqv1ucebIaf9AncpoABAbwR2KSjB6SbKVM
q29W/3ZLBsksRhRM19rvkvo46AO/vzjqz322O4i+xBPS7Vd4d0K/2ManeHzSY6oacU04YXRiuKa0
iNFoEqKprnvS1lVLWkIRLZrPXxuhdho9KWkx1QNH6/7oYN8C0ECZDijri/LloZ178cGLHxMemDsk
hQuuyEh2ZTYerAU9KTDA6wCGp18tH+dSFR+a/lVFWcRCeq3ov3h1otYui6wEmtLzJvhsmD/CmmW3
Wbi629O/hRepWHUyUIXlB6+VJafIoCTgBXf8mALNDp7X0GHVD38s7OwzZZ+watBJ0sOgVlfomPJV
DlKCBIm81KRXq6MHrue7Qz9CXubToo9xUBjB9164wtj7icKKih+CSomegNxQ2d+P4FBjc2Mmqm/8
4fuqI3tc7Mqu3pP9wA/tP82Ty2C081iQScWrl08/nHc4ipZ8HMHhV+VJO6vqOgbNlfKZ/3vLqYbR
XTZPbf1PfxH2AmIttw6s4J3IurEOj7vAqfn+PsZlILSWgEFwI6ZzZOt9kE5bK/BzQORsix3ydy44
ldrlB7rnoX64UN3zLWR9LfTvQLyJbUZWXHGMbeP0KIAEVWy+n3iNxhY+lfvEnIBNbqCTVtaj4JHJ
tVUNvD0jwBqsyv+lZ3bJl9u5N4zCFx9LsMpzvC+GfzUzolG0AF5RymVNiWFn/06hSvsv3ZNYRUuR
5goK1g/7RqBdGnV6pT42MNZcHZeCRifsFIkSmBLYTkSreiqNdQBeME6j21VgkIsXQ+wJAwRdjgFF
13RzFy8kcJ9+oXLMPiv3bNYiEO5l0G5N5eMpO2Y/oO0LhOyCbODEwnadz90zisXM4tkdN79gYAFy
VjVQ5OAchcW3i5rv5j6N5RHZtrd2WP5wXcKlOKxoVa4iQ3EK8UnN0O9jpd0FoEh4YlmGrqYyF4vF
JVbvM/Smu+kdydAfpUBK+bj6B6OeRoNkbuSEcEbLhRzx6QP7Y/HMJu43SuKAcfqBPGzghuSGV3Tx
HffKJi6jqpAOTgTtgcBiwf52gxQ1zUDxFkf0UWU8G2jB1oVO2K2lGqhr3kFmbTS7NKnbjQfRXCLD
h3vLVZkO6jOr6Az+sxuzywF38rKsfqjzaG/9osCAuR4T47uCuQB2cG3tni795zQFDojsMWRs0pS/
bj5v1t+S4xYKZmYEa1GsrevBUcIRQksZQjL9MRUJXq838IKZMLl176YfmVgt+qfSzLY8XOZ1Z1Sy
rG06fGG5Yhs8UIrfILUY//tRsaf/FrBH0eDhnQ8E6nbdNMcdeC+W/VinNIT2X1eFE+B2/yue3/7x
MfUdOC7KJHl2MkhCBztWw2ogOcoa5lgVSklfrr8jO2QiHGxffUhu7vgOxtsvxna6BtAX1zZDBmUV
2OdR9uq/GghEqRJG1A2y8ycc5FpbNmNE7wrkp9tsUJU/1pE0d0Kmdbj1x1/FbedGjuNvgAN09Pss
Kbh0Qua0Z8i4t/ESX+Lzj0yBz1hC30B2jqFYzQHoA+nK9re0Zs6tzNSzZ25btvG3rrGkDJQB0mUZ
SenOmLVQbhfu8ddvDSSbymiAXdWPBWvBUU/1TkcJAF7b6DA3uQVAeWVSsyXZjT+/egw8xKSC7EcP
ccIpV380HcKRbJw6tiCCujUGwDTrraL2MuqQxzOWjzdsvjm08BDxP705b08kaXblE9CUXd+kp/t+
JwhO4+4SKJgUPZsumjVY5J20P64UNmXn+hEkBU6lBTOu5btocG+52B1/26vI1mGDEU9+9jf/XzXT
T48LuI345s2Zkbz/Bk5JIBmHziyiYCPsxVu0dKMNkvFtQ1M7fzQIjlT4bXbUbX/HTJbL/M8TdvlZ
7IDpY2OgQ/WtbqaiG+6MK4iqplbyXPzE+X3NJLjQ1sWZSinzPD0XlSpfGUL1ht7jGP50fq59VgY4
3HP8MAp4gExBvgTOuP0w6Lpm5JUSHSMmjFbT/cUMBAuy1TMpSWoTKQvPS9ErFF7Y8XAgs9d8DBxV
dSYPOOn1dVEITpkiCMEdENdJ+BgdUcJjobEscy+raxy820ddWGoKDAdxoKIkkddk7m3WfvjvOthl
hDhh6BhHzq6weVSuz+l/6tlmAdJrSiVWog5FYoonemA5udxEzeaFrDWBi/T2Xxc1XhDV6hZv0kJp
0gTSqaDQB4h/EjaDp+7cFGzzogf3NZmL6sSyLv0dNvaZ3iRDtw6wTsBqfSZ7SDNgQqKxlmbiyeVi
S4ltNodr58WT66g5PwQffQ0CgPGNu5pqYfVubDFYbkeMECJpviIszo94b8VXP4TeRkGrkbwcS3kk
39SBTxqFnbQrbcWEwwuwrb0h5cFemS6u8cPZTTFtKdFX/9P3/HBEfOKzDLDH5VW2lxu+ZgJ5KHCY
Fv2G1QH7w1oXV3lhULSgER1EA1128mKUU9V87OKD4PzFxLFGNv1FfA0EOholZJbmAvEHDeiox1I+
WexEc7uZE3+h+cbtTjTT0vllXLPaQR0c3ftU9r8HEEBZGOi2QTX8dmC9ybftLpR0DvEw6luzVIfr
v8zneJ9TmEQ6MMT2onFrP1siKm5/rYHOY6uUS355Z9npq7SFAj1vwkfz7DxKV8cb5A6vS50n56Xa
EYF0HtYmUfX4gLFgWRwXv2wLyAntggcSyC6vU5JDDEIrdW3b55hzGNHN3bPhjO5VacpjTDbb4rzT
RaNNL1HYy9+Y3tdz7hBbEekeUYW9kgBsmXHGiPDA9EGx+vTzUoVIu2ZKA6XYq1VVvmB/6J3IETfM
jziVjYSHEAlDla0UvgUozjfRDE+iv0Q6Tc9CfWBjVDdOPDOPGD4DqGgkVr+5jxVHVpI2N8jHV8WQ
N7uy61ODG+dq6i7aChuBQ2cyaedBwF0AoChMkpkve2EpNJ97IIp7/oo2G8zLgRQcbVIb/zox6B7A
oxplR2M0ai3hsvPE4BVNDNrds9JmyUgKYNc69QP0pIIiLCq6F815aK6mXYe2R6+WmtC5zcwt+uSd
kJje2Er1Nm4HDwgJaZnYoGYMKEkLXESLyvT7S7wMefMdh60TMTcaeYA6otcrK9N6ca18ek0zbC3V
OK4o9rRkYRvZsDedLQfDR/b8zSkez6hoAX7I59LLi0Ua/6P7rRdrAn9DsflPcqHkxJXwRbCGkkgV
7PiY2aoAktHZ/fLZupt+6rc7B0a7f0vo+9GxOMXfuVChfuFz/yyiAjz46ACXbLN93+EGjxE7kUPE
pn8PcCH8SfwdZTHpEW4in3Ay/cIvco289W1E5948WmA9aV6YO73Z9wVu+TpvbdeTFGGV4yl9qUvr
yudOVuP4usCIv/9bUkRWi9xDD4umKaWrBhRQy6dP3DsCjeAPXy2ksaNNWjVtqyTS06VYd9YcEf1w
eU201SLY3SR1Xh7UIK5AeODdGS66scOIiNzUC8MmMm/0RIaWfOSkDa82AXAj9b2V7t0ajeZZnQN7
IyoeGazrMlrJrvbPfOD70l1LRa5I9YLU4EU43btmOLuzFGIbCwzGq6APu9xN2UfJzJK5NTEzXO4f
RjMh1zXTCPTOoOacpQb/A+6Lq3J5XbqSI8OI4m+ZEFLQi4YDFPq30uKjNLnLjP1TZliFMIbfuwPh
J6zSo5TdcXu7DTGqbJDnAIi6a02/qqr09WPDwnFdH81m9uDqaN8XhjRg1iKajvsgb20gx54tCXNr
l5AZN9AFz2IFMDz5aFr635m9d15KHHW4yERpEAjTG4paXzFWIETyQG43fQg0mNOESsHFqPtNyKb3
zQ0Eeg/Gp0HDozLo7WOAIxXryogIWE7YFqdtbm0S1P4diGZ8kAlX2psYLmJzDfGIj0UtCWYueWY/
4+JwtJgUhpQGV5Ipaj+WYB3iUQ6Qeqb6NP18D3O8rsChjCG1LW99OOcKAPY0jLNgwLzmcAFZDvaO
Py0dPQo63YRUTs7bXk4ipZT0w/Y8IVdVyRRpuSWJhAn9KqwvnpfNTKDgNjptF5OZiyCmBjgYXEGD
Qphe67/jv0KLZT3BK8Dsm65KG/fR+xSXbKKd8jAk6TcgahjMBo9mf1vy/paSl2FtKlSgyMVAn7Tk
bYWTOZLeyekr289naU8h/Rky+ZhcMLIJpr0E4kQilA3gjDPBquKUqvZQbZGHVd+cFVt1Wv8xBFZP
UqhQarM67gF9tKSXJRZOh0bUORWDtRz7Tu/mLVNcgHkeLJT+rqfQJ3urzvp2r+1Cfzd5xFHdn1TC
vuJxss5HlG0HWCKN4WPB5ixXyjmirEinktZWqmBGCigNwqiVkR6jX79rLDVUW/R6U7Yg7oC3SWOO
Sopvzre5b9CUd+klzjGFL6Xgfo+7pizz+9wOe7bUZqDzFoiEG3DX84uHI34llbOaw8b0JUhZUFle
67dGNGZ06ti1S2REkFRSAiYP8z3hPoPIgT+lrbxu7tRDjlC+GbIYnVbU64EnaTyHpWifXuk6Sn2D
hGDYqxqOeIESLqdOlC7yqgisugDK3NVoZ/gSL9L6nyk9XkkSKvhIzoZWaPb6QGJofxgJJ3mP9M4i
agN16GO3xBroqwjREWYGSMbKwTdJIfsFNNyqWDWBFkzNvnKnRyBhDUZFIlU7a+HmGcwcw5fIwAtb
kHZdM30FtlbXZhEDCVF877vYU3kDX1PeUEa5uuAcu0whDiqRs2BROS0vJFPVA6yuwB4eGZWB7RHx
GLjMREXb7d2zjVTqVptu0DWajMyR4w4fgRDRFkIdhtqW5ahgh/Nff4kYJq9OsGejhm6UG3GVqwn5
woTdH6Q67Yyn5C1upnMlN4m64lUtj75LgBbdwe4Xv2VxrhMP0j1z6nbF0qUK/bDQ525XEsHRclgS
b0iCAvSOoc6HZxeMArNnPZg5quBhDhYYSpDpzZ4L+qMdy7bnKD72FrXywDDyvDp9K7mfsItlRL5n
2Inu0wxYTsMpYC7xAjzLHWhMIZr81z4sdXD9NzMs+2jojyQ1/mpdVasFgFRTGnM1eWB67A5iSo3c
Sj6GqcniWeOixW82w8UrBPkb7aGgMtYvTK6rIOfQcfVWLEFI5mGVlTVtDPCwA6Ytl786644Te0SU
ebaE2vi0a4zyUXVKo1TJUFpJEr0Y2ViwUD9WEJdLYfEJtN2g/IyyE17jAFF6cQfmLn8iw2g2TVIN
HbIfB2O5vd2++D+Ry6UbyyK51OVO0FNbdJeDOa5WmQtTaDXzisSr4Bqo8kpNdySQqd1MewuVvWiG
QHmv2jkpMwEfzlViHBogSbLb/VhFic4gITcnxz6i6Whqsc6pffIyyx4PMFzTYRBqnUxdVKbpuGrz
55F9Ephtz/HPbONhSJiqnIjuFo51DFXBNdR0PRJwnbCj7FFlq8ESTWMmAue4JCP9IMCkjQ5MOMgi
axXnT6aSfs7yenqfiabdTmjTe4dMrvr05O4CqkIGQabO74GODRbJoirr2uYYHWtmWCMZOkSJvezA
FFeo5EgF/PjH5esE49UwAL5sjVEcJPf7Z+cwl5uL2zI3k/008hL47o5n0OomwBNZhsC6NF6sa4HW
l27XWG2dtDQg4ZjGb15Obtir4X1ehyF8xsKdbAD49idKLRgeS+pykv6+rLQAVlSnN6dGCipVWSVW
xvXqqEY0waYUD25VBuEPf7CHvKdZTnC5w1jrbTnx3TSxhDEKNJOm6PImCKzWA+qEgfse1OFARP/0
qgFIzwOloN38MxXWQzgRH0PNp5QBe2KCThI1wxSPJ98xERqBQ6/10wc0ahvivHUF/dinzJUHhCkK
pFmHVFbFSboLwNNi0cQFDKQae+iRMiagRxih+54LdON132PF4d7iWHmkHxZeyd7aH5F4xfyFoin6
9xMuCgaYxACj52qn6Is/QulxmlN4ejXZfBHElmwbgLLofxJNAMSnpT+feLoxTvEMD0++sR7HtTES
Sw0y8DrzbWbtxucRsXJ1oOsuOUM+tk6H+uwoC77z5/N1DblrbU7S0dGjqNrJrM8fozJ40Yh9Zl4c
ckL0oGaFPRWXAyTEfR1ra/AVwSl3MX+d0SynUxDGFo+Kmz8xzGTRyAJm48jv/8Bdz/iN5BZ38fmL
s6qy2ij3y0Q9q1RPPXu/S1VaxZrL7Z3gpn3D8sr4yVGlUcM9CCmd2GZ8GTrfnFrdL1/RI4aiSMMV
/Bd/FfwagP3jMcGkPCKmlXBXtAozD1ZSisbUUOdoj+6e8j6yglEZHf8Pmt1G7hwSMxe3IdSCKCYq
enYz96tPWWVOUFxwId9Xzr9LnDy6kSFs9tuBAG6Hg66rKOvlWuCqOC/2voqFj8nk9G3m976o3FA5
dDXfmIomIIxaO5IcfSU+7WHb5KhcHZbMIK0GK+Nf1YJsabTdXsa0/AUt3ab8TZE7oE3WGFqsIc1n
jqXNDvEKJHH+I0YuYXTQF2Z9S13TniAGu9xJ7zM17p4LlFhKQ7pAGQDJM1lX4UahxWQFcKgeB01w
GvtYDdzQRWy3kA5NsCJfPyC0cLEJC3gNm0SfYHC+bv9Dd+eZUlvHMyj+6Y6CUhKqX5r4Ea0RWwzi
6w01WNpHj1D1JCV0q5sCroBBNKJSB/2VAKj9
`protect end_protected

