

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SnF6N5xaPbBd3zdyLJCTe5J3pbcy5MtLlV0mA+szPwmOne+iuDA+SCWteU2EEZDIYrB9mWb9yR8q
0AKAHpZPGA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
haVc8wzStzlg1qKktcHL156SRFqTRBKPce/boX0HKziie52LAZdHseY5z/N6Cc0oLr2ZJbzqSeEm
+zeAJz9WV0YTI2qvVbMq4XUBk5OpmpKdb3ZdliVlfScbCKhoZrfQdCAL1RchqtRt1UZ5NTbxPcnF
p5aze/h1uePyc/nImjE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HbOt/yK9abjBylOCu38tcAz4BNy/weqeg+aFXYu8NPFHmPz4jpKJ4yoC/cKNA4fGlORBxz+FO/g9
8Z8YUOaUR1cq0M3LoUZ2aNxMRjv01hi3OMe/zKkZdKrnjQgg2t+vAlkxK8neGN+eERwXRqCJP3lj
7wiKWHik5U+mspdaqKON4/soRJ623Vp/H0Y7LmOLf/UodNxUwSFNFhQuFyQHHwRfbiX5oHoGfVJX
GHJ4Oot4alViRR+a3cv/wcjJuJ20V3p31WM6PpKjioC3YqrzEXxkwMevbZz7pQBe+t+T6GqSXt1S
/p29OAYjS0qlL/uqmybKxPIhSr79b5Bv01HRKA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EEAnObxcVE8mih2cQUC2xFbX5KRSOdfukckJbjcRGbVu07Bfpu32rpUwfbbHUlwDpkwnrbwMaUGr
EiT8Uc1MHbVGHcr52UIGwx1sJ3JS1uBrihh2ptmQc8LQ90RGk5xq3VE7apJjPeJuwSbzcIT0IZI2
6Li/UKougJYm5IEZcwTJwSceGZFZsvdEegHRlqk8wCuepckni/Ttu8QkXs9mfIcaKkcyPSjlFE5b
jaqqxp7rt/QVbzmsRYTYUe71DiiV9B2O+QHN1ksLsw0azMoeZaluU2e1kNd9EaU9T69ahyPF6D4U
N8ModewQv+LgP1JVIQdJUzHuoo3eN/GW+qDvpQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UAjXKWDYG0Qghtr3vhgiUwYvolJGnk2RlGmS6EIXQrOI5jxgSgdrrG+bfBG5EAJo9Hp0QOmtgBO5
U/5XOkC2rF3uHDSENIp54t6Q4kDhgvm4WMOMKakaI3N3TgMjjq/0xinfB4HKbc7fWvsNBmQ63Zmq
puZ0YrBvXLQpkOZfblCMp+gpwyrQcHJQrUROfMUH83l922y3MJ2gfMAm3KZbTaSpdrdWiOvvMoV+
Ze3ydpw1pyQE0xf476c5LlrckNCl8ZEE8ewdNJNPLwMxGo2gEHAU3YqkkP7puSd4zM/mslX02xXA
DWaa2VMci5PGyNBJRWH+i5ZQpEHogv0lDei5eg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j3dzWgjwmtwO1dLyLTvf+/1Cm8rEjNLd3T8f+2xXwaJ05VhftMV/cMp+NFceRD1wM4+ljPcoxMMC
OR9WojcIAp1NtPqmrumc/7l2XRjn3rV83SgJbrM+AjgDWl9433MM9nkp14RfvlTxqqSRLgkF3n/r
C2k5SwIQ3TJY2OucIq4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QmCUZnNERmx4Wdvy7fUGELgpyCDsfRwgkxM6vnznQKlMAbGk2Porujld54m9bDNLddKmnbiJetIU
KgoH/5SDtatessfc55K4Ire9g1rDNu68Ffz1JxGatl9AEuQBI86sp1xVgjdrhJVNLO0/5/3sRYe6
MNIpy3fVuFR5ta6FaoJPohjYV26JmQeeYUvZkbv+b1oFm9fFkS4wW86uqcM0IAWWmAnEL471AycK
Vm/Xhecn4F0LquXNL7Vy9zL5Ao6YBUQL6MXy/hQ6WEJnrsOpqMI27b7XQGvCtPzK6Grxpta8cchY
f/pyjTZLBinxKJYzF/8LUSgm2hpij++e4Ty8Kw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 333776)
`protect data_block
y21lc28oMEHlx7O9ax/dwdpcIrMu7mdyEuEzeXcUg2FYmLgbRMvGYTPjaxAfUysuUoUhb1AyV+AX
vUJltWAEFmKwlWnBZsf5lUrzdUynxbUPHKnDhvFXAWiW0ANC/+bHFJeAOkotWQgIPPcQyfKWliT6
xgHMWuBvYw7Z7mY0HrZVqtZjRDA7OWf+TB2pJaH13bdTFko0/1BrJInG7ou4rn7i/z0xCKv0Kdfa
jdZyQAlvENJmrYUTjA0lYWQsO2LH0V598Gba+5FnHby2RgnP15stNTnhpUkSE8bK60r5XEZC+ef4
4LAF6uP1ku9Ei4E5dlc1DSV3ZNfKUKUZr5LUzmDnGR+TUAbn1Ov018V0S0TXjwllCPo+lJi0n/P7
F48jEmIOTSh4E0HSYSqdWnG5H1298zjOnsd1CRpCCerxq3zOFYd2AmeFWpAytG6Z6QHNfq7XI1tc
CHeVcTVOtF0sjSQjyybymNWkQFwjDO5ghMOrOAiuntVLgQ55Dl2oFZkkc+6n9dMOTXigL2Xm+YX4
A24CNa7/32VNW+O3tiEnLWv1DBI+XxGrheBg8qkJPCDsmlS+V3iSLsPKAClRgDvGlJF1z8OaNi1q
kKnuA4m81iGsj8+4tpRTNyvLE9bg7agYDIW1yUua3t9rp77YLF4eWaaFTZ2QySR2448N6yyN4X4g
8Med/cV1PtL1ygEU9vPMcQDfZGV4ztMb1pMsi2CgK1ebzUZpdmv5+om4BRiwGPmdkI+1dP+qieSN
z84kWKgN4YMHn6unq8+DVtY30R9CvsZVNNBN5qFrRiJdDFmhJ54v7GS3711D4k4JXWkFIXOjwz21
11a4gDQbHtBve11TRc/lJv5LfdWG47TiwYHRY/fHyMWII/9yceOqwZF/0R8kS9V9lOla1QEU7+K+
1jFVwsEVbRtd+imSds+qAjOd5/0+8dYWP+GkA/NeD6/mGmWiE4m4FASMHFcFyPSJJECTRmfMRRBJ
VdV0EvpPkzsFbm4ZeMwDalCz7lEtpdHs2/Ixpa53US6f1a2v94p36eryiAR/x/yf7SPDH8BIyjgc
SJlCMYMgnMMYZbi/5zDoRJCfbWOday0tVu6ZRhJLhPRReHSAAodghUPu1jlbKt0utweYn8Xt87Ln
bEZ2P9mrwDXUrWugeNy7h86QdLKt5TGMxge0qMPYzKWPhdOeGYzVcqtEYUoHLnnWvpUUtiO8NPMS
QIB4OZ3op6r2PDItxt7xacYIrfPzloCV2LfwtbinjVKl8NCEbi/T30mu7t2d8vhh1QmYTZzgnHFb
sBNSqelILQfM2GUR3qfAs5uS5fgbo13SRBGz7W3OpcyrhAXjNWshbcJNEhL6j8Mf6kIgEzN12rUb
dSBFhl1NLNHpPWLkX5LvbeVZQUfDaO+ZaLKNre38U9y60MBuY2O44zLOA5FfyuNqeIQyZE8Rcs1g
2nD0YZP0iIWbJysSvZlQcPQRjhJkiXCSerh1NDcT8BYhPThKg7wFlH3/E2g0XmR/Sq/pmwPWcckT
x58cUWmQVXrkjdTWcJT55/gUw/47axfwn0TkgWwAIRTUZEed8k40YhhTxpu4ekh6iPGzkfbTFJGC
PhznJjpM4dLYx1bdMy5EWavTQ35A2lhOKBEWeOZSkXeD9FNkIwV2XLNnDtjuLR9nqkxGlNMQQLtf
rLGrBLKKCBNMniMy9wiSknpmwLXFpTUTbDxTfNPQpIDCWoJKfFnnmfJcao9N0pXCKeg/9K2Bq4vG
ZgOpDJAMbl4GSlUHjSl/fUOxeMZ2sfqql0ZWKqAgHkiHfLtA4iytlg03+BWqIOggjhfe7DE+zf3Y
LBXqE8cj2xePz7emifk3C6fphb8KfxVocRH8GoeQYQ7P1hQfekELK1TjSnslC8xcbVNWS3SKdjIj
Ujv+oBBfGYEcA8W6s4Ckb5WYuwSwsVp+2BEqDwdEqj3qUopiTOfgZE0idVsKrxIPL9MjovHmq8VP
C4hxR86da1jGi7pcLLRgaJLiPbtQdhQOmoATglcAgUjUqfJtRMkzStA50YSU/PjySsvkyDvv/KC7
8/G0q562pzw9b3CD9/SxNU69vGKA8Y14RM3A+T15R49RlJwnYmGRXWl+jQ7xK61fz6BbvqCwEQdJ
pir7O7cygt0MP8HT6yT6pHhS2+qW4fH4I2Wv3RKtVoJMARtwP2yYjWwDs60u0auWI10XF3/wKss1
8Imw93Mr4OuHMINs8LTKZ0zwsEaGGK5UHSqeENlvQONOPcfEq/dwPcStirFYbDYpzXEvLAjF1teZ
LNbIsL40BrEmpOWz0AzajYrWQ1fU/cZ1EhYwL8D60U02Zygl19nqvSS3ULnrNlqduDLK19nTqmEi
84+1LjTm86Skf+u4efnYjOWRZET2SVCh9SjjgnYx9xvK+SQyRzyf5UeVZxk4UDAu5KA77bDhGTpp
pnCLc6aDb0TELlyvLXswupsqMbaCUys77edmxMoUzHq/8Bl2GB5582ca/BlnYz7DCqbEwUvg1v1D
2RGpNqmLnH7kIuDrwGydP2V6SHXYvXxnJU0i2ScKDzFraov8DE6+aqrctzMMjBvTvGjDbDXY7Kz8
BJVFRm6/r0PwspVXZr/oYDwnVQ/Qvlw+MolR9xRIKgYI0Uxhijy64nVBXfc/H247argimEAxbTVT
OYYLV1vhBZg+Gjxqadts7xoJ0g+X9q4753ar9ynI4vFQd9Xfu9cOMAuaTZKJpeaG74SJ37z9kooc
0zKIa+Ae6O1ZUVwFSkxYeesJCWFlOiWM1xrjMUuqS5jGq1hQMULoQQUeueHsnZjk26Kkw/eZgUiP
Ny532prO5eFH1D9ViKS5VyBouXASPgRuYAf7D+hjNT0rtJgCuTlYgmMwOI6NFuZGrb+bWtcIL6RR
VFzo3q1x55cay9FlRcefgrbl/vQsF+3WAY4KQ/iOea6Z74xaBHW7CSpXsncyJrDZ5S5q4HwdLjgS
AbhrEe62p9b2AwutpcY8KbnPdRFrj9OsGw+1LhQb5Rc8FCFxnCBtHpVlVKu0ZprKyUGvRFyRoVof
AZgsD2HF6ibFS88Cp98igMaE+zUEaaMsyCu5co1QYZnNbp+Yzmkzrb3V8fCSC0FdW9H7v+SEFkif
24rp80qsT/7oyCnzF7J3jX8jkGr+hR7ZmPufCHuQcPuvlLp7Gn94nYM5tMQqSy/0csFPjegmKJ43
gGGTbZkr9bg+bO+ZGI2nQnhZSAmsZZPsrWSOVDNvcqzZfrlvO4yKVbCa6xrYExhEppqVZviqkIFd
vY8oHIgwjJfVNMu+7z4aH2zLjl5iXCl5Zv8XDf8Gn5bCVl8yVGeR9Cw/9yke6R125tXaw+jrEWZX
xSe/ZGvfWNH6FPvG9QmeQOX8+E3DPwqxk2fyaLZnOlmuqMzAs4dtzEhxBTMaqnEHa83zt3Bj2KyV
OyrVkcXzTErza9VUjhzeSbqq1b79qqHn3QlvyE3CWWxkcymmBp7d4Qi01hUtKhl77ZAW4EqsoUVb
gfghjmVFgxpw5hWNfEI0+lBjh0zE9AB4rXDy/b8Qcfd4ra/0rTmHrOL3ZJ6Bri1+NzpmmVVDgnfb
UxzVrDbqQpbBm6r/uh0NaLIGlMqqlHm4UtDXNNVioACoapzvuHT3bM5ErcUQLnogaIUpRTRbLG8W
XqWfo7p/OzwITAFZO76Uj/ComA6uleFtrL7naAOPxu5yAnRgsBaxNRrLNSN/Dvath9pfFMZ/3bAk
z/WC5T+HRl27uasC8Vdu+7+H1fHO3Cky6c9NjSeHgrEq0X0MlMqK9nhf/7DbAAA4DLgI0Ymy58fj
ZWokrf8Yl5x5yf0KvkqiepDH7Olo9dZgUHG5nCHor2zahFLnNBvQqHN7mVwX1N3mL8iex40c4gjC
zi7W603OzPElIhW9FyCmg1+Q+ht9EZqzX+zo0Y0DmIw5vSIqJzyyQ/ecd/qFfBdu17u8QxvtyGkw
z6vlwtIBugC+3CUsAfP2INjf+Mh1NGoN/zFmom1NoSnCaDldMuFHGkjgERgVCPP0fX1luUhGNOTx
gi/p3cAtLHWoIBpi9LS3nf+qCwxqhCsfwhuELSJA7DYXuwnIolUdk86wzSLU/JUGsuIDebvicZ2E
e+4PYZNq8MTGH3jRqwBPKVJo/GlJGMrO/4DZr5sU809EaNoPiI1aweJba9vbsp1CP1bP4lAwxBUJ
vWwqcnB8Y4chpNQsRVWoCadOjFmyjod8I6Xktmm8w+Vxb458d7WzIMWrZSX2MxH4uc4gef2Gb90L
PYL99uegYeihdwikTSg2WUd7ou0qqGpZrj9e14Y89WVheiT3l7IlJaCEanK4Nvq7YawlKHzF5YcK
gSsh44FFY/FZEzUHZsXfPujL7eh9fW1jazwlM82GYVeNlbuWGEowRzr96WXoAJfbw3ntCyosFILm
gykc94nS9Ij+RnUwdY6XHSOdG3vki97HG2Rah8iCayXr/SwCZyUWtU4ieL9mL+FQdzGnVOdOrsuy
SPL6mVkQwfCTyTQEsVh46RxrV+cgWeLuSbAHuZU/alb+h594c6kJIQ/uzA3lpRKFENTJuIBMsN7j
Gfp35ucx1A9hBukIKh9e/irL2XXMU/80dN65dh8f9dkMPak/V3SoD2wCAYJjYhFAbLWWTazn2kFK
uYyXABir4Ba/yIMEfMnj3NW/sdxSmizeBGeHdbg5tXa7p9hkkDO9zfSWJRunSYj+avGsSRHd5YkW
0onDgxLgzaBquv5nEcF4QLz0J1selVdcp12I3c7wO3NlsebxXquK2Q+WAPurImptdqWAFIXSQW9T
0Fs93fj2VsJtRqDuR6MHEMJyL9ORRSpkPC69eWRgbroKCzRFBbwSDZWJ1xTYdhvP62PLyAhzsCah
IbDaUOEKH0cka1Q4pekH6oKF5iNmPPANxVhhsPhL4ylrJieFvX0LEF2OHMI2Nymfj787WcnDEFyl
r0qcPLIKkVeGro+P/83bxUmskTtBJUKYvBZuRQKKOyng0Hz6Xt1pwcTZnZgPyXF40LkGeOJoFxWb
sqUtTdHTwy9uWr0Nv758+GLapvoHtZgpYHvNcMSsNV2nrSNb8P2/Dk9nJyGEGQYc2HlCToe/TadQ
QQccQLZQ2buyXODj/IeGA35JWIz96xLigH4k9aXenXrPW+9bX20M8FXnqWN/FvC9GusvgxMfcOET
664EyfvWaEmxAq9X/2Th+A7O7NsRtz+Lz7ZJ40Y6uQDxpXvMU7j4c+dSc8zlfZGnpMgTR/cqgKOl
ZPdpOrhBl4ohf7OzBqjehBuF4yKIgP3ZjOAq0KtFNSb5FkvyvDIwx5spNdLRx/gVzdjFNbArC3zm
wX9TQ8+ivBTWSWXuIK1AjBXG4/z6D9BHmT2B9xhdJigsqrD3PE9X25sRK23Q+W2PMl0Oy26DbyQh
1UcA+y9vIaKVz0Hf7YIrQio8h0cxdhajVHSmez2wrmM3xCa0e5cEctjF+wyhG4tcpc+ZJjn4weDe
g3TExpW0Faf4ITnAZGVsaGLUH4FIvupd0zf1R9Q2yrxOvOjCm8r0pZc6FvD10xIEpoyBaxyIDs1c
j3H0wrQbFaYb1Sf+tCQQIJA8K69gEMr4nLURqfhwy4vyquXnHbsfxCDjojIS8VVMMsvQ0j0sHvBe
YbyqDA6ZXfCuRCsN7frz62VO/LQ0bUa5rp3gDNcr/X3ILTRwRDT7kCVPAgXspMIeSYCzUmM6Ygy7
c5+nvX6R/Nm62zhxJO1wpphknDcD1tSl+eNVh84omTK0xCLaMWc3SuC6eRc3wlN4/jaJnlzhgpOO
wBtYkwPIs4hj++VUCjEaYndtPXzrei3PMliXoeIUV1l8fwD9hTgsxiMQvBHQWaKXyQ1jOl9OB8gU
D82Mo4+F5i3dI8Hlfy/tdd/wbKd8hAMVInyHRWqbL7V+XWMtddkUYlO4VTMqn+ARcrzlDr135QR7
M3iMb4grE+DJzr7/HBp+MTTkEBF5RcHB/7zA6JY9rEz96AYV2ZwEkr8436kvZVU7hahiVW9m25en
zQJSICxNom4iRZMtdGsByEilYU6xzZ4JOcgWd+eZdhVcR7YkHW5CL2pXptRdcSA061pnTxdhjlqP
8gMEDqRWxbdIHArqoxrvfgKMVFkKL5CgROb+/bH6TeigxNSvqGDQ40l81HASYfNvBG80gZK0MiD4
cJ/BKmgIPWIhWVpnRklpvBc5x4yQV6cUvWmNn55FEknf0qWzuSjLLOCaDkP3GYf6K/JOGG6AlIot
lSmHhB0NMboWOXLdMc8UXjNbZiPtB5TRjrd2FNFyBQYkoYmtWra4ew27BrpvHTuc+zTz0kcRhq19
7aI1hNxPl2y1w9KaiZLL4DgD5mbAi5JixFrMAW39SZslNtrQXqz1KX/JGoaDVZG9aVXnOrhN3qqo
kj9bEr9yZS3OzcsE7dvLU6AMn0fHmV9yXLKz6/7BDJsnwNOvafePllLxMCboub6NOB0l6lgXLuRs
RuVVIbLzVOkoGGI3ZHqanqL0BvuITtNZXZSJNgRet5KooUBnlV31kTy8/Vys9xcRCU9apncI0Ca6
GA+YIjGnIUFiHr9qwTYy+M8LgpvJ+5QWNCvkaV+WQSHqJX89uetz6MjQB4mkzsacAN0QTvox9ZrJ
IG+j8pQHQU3OUi49ii+ue70HbwC4EtKc83UxNOVhW9AZQY+D8X1HdvCx7txEx9QuynyaM30ObpQP
Q0TorY+pB3C0yBo65wPqnc06jPcqTKI3yNOqnd5hvQjgltBA/p9TqNiOAQG8MajIxy7pbAazkOGV
mDt0CRMhqi6sXF+70DSVM/uWl+bwi44ElajNKNL5PJTsDRc9dleLsmwjGO1sdDbtkd9Xuhye0o+p
GxI9nDa5DqBpS9YtdbemhKZMzjEr1RlLg+f1g3iidFBU6YUVRnYqj5fS1eXib3EpE1jludduxnYB
YMpiHFs+nUk4QU3qvWxNh+IwlypWvC6tKCxgA5HcZnW1gbBHmzGv/jlYGxGKyl3eiGW5yct5yySC
9Lb261nMIQJheToeWBOoQKsYVcATc2tXQWp/fGvIFHdfGxc0GVS3l9/GD94wF6V54Mp/YQJdUb5/
vy6rl75xwKZzNAU9TKecUZq9k8NO8O0VPMqwMk4R/WbJp6jjEHgCvd+iOQHUnQu2frY0HMd+2Cpo
/GsNU/2fqpxgBtcZIvJfvc+xQ3QPLxQaR3G+k3khddz5dqSYRkHqhd+uTWWCM1R158yRF3AtErYb
PQTBiLbonDCcubxPQI0C0+gLjFC4ORU4QLTMqtk/U0vQ9dMwniGymr4Iasjye8LL+2Y/hDP5YD9N
uO1X1fuHA9gQw1ppiL45hBlOMgK3oUoFjYx3Gb8xjuJHM7+zPa0aIU376gP/u0DR3ryXXz/fr2Jg
ylknRwGAKl6smvKJhd+/pTKCM4Cc7OLOYUNN7f9E9pEHFkR17lDqyiZRkrHkBbQBbDK3OEY+rg3U
jfXBk6wXtlOza1JDNV2jO1y6rF7z3YL0uSpUkJg0duBACsfDI1dHtqT0NN9nHP11dtjnu0c5/fai
R4DRosmHj/r2MTdUxTVrnfy0sQvg7B5nb8Z8Dz7dzpHuH3Gjf/OA/TO+7NQkGNZcq88N1zGfA42h
4QTzOBlOaFP5NF/BynUusO0dX8YLdWw4Cum3hi1qN9VWLmwI9wk/FTXp7xSxd++4q7TPAvc1d6S5
ebbaHPrwTm8niyJa7tu7uSCFEhTGRcoWa5AgxiA/o02xJunUoraYoO83xXM/8FAAjXOdiku3Qviz
g1Xak3ChhPwCr3f02uM+XTH+8VJToYAQtYWaqG+KplfOCIG+oezHuA5VV+n4cXLosMViwhtS+3RK
dt+JcFS/Yfognkv86Rw4TdjeXk+cAn6NUVwpPmepTjYALT1uI4HOWp+dyTuE0P2M+TbzpAR+L7Cu
oJLGdfNO9CuJ6WSKMapKY2zfkLtGcYDd6x3S4UBAOAbPHaGPjN368+SQvBJwZuU6N4KPWVLaOosJ
Ajajvo1S3gc4S95ctTaxnCrfFNy+9wtWBnakcD6mM4KTEK06mI9KTUzf0GFnrBuoBmFACcTJSuV0
Q6tI95gkkjLvlKrFc41ld+MOjfj5udxDx15cUX1L1HiNsMaUD62JMzJ5YfqihCmrnCO4Adr6nJ3p
7GBWqrpm3NUkQOnB0kXxNxWcXRaEC/kdhZIbmQNcLTsAHOY31ZLZ+6lZFheFNMVh7JWwB4FHrvev
+WpjNpHla/UiLg6ujVHmHV7OgJifqNAAquI3dQNAHyV2M/EHTreg8QVrw/BcJ6NQhQd3qqoYbtWi
FeNMd3CLlBr4tHclGvlmQHMHXjQ87kU4fANMVkza7ix94NU/hZ66c8Q7iLraSk4gBDyGKejRZ9VO
6bw5RqGUlgWrzm2H9NhqtPq99CLEOEpEC+ntjWhXxMva/6Ybp8MwAeRZFELIjNxcDNnEa6Z7lOoV
zaMT10qx+7vyC0P5BbpFeaE5cNJI5P6U486U2P7p/IQE92Ms177pevu8/B1L+b7dbk6mtNnTeWRS
dxHo2emCNHdWjAPdkrmQQ7cnKiuWuZN6lEYs5eUrhxu+qWMnI5S8kVQibvpvljtgPOBLmMwqJpHN
cs8KyPX0omlI7eYrdXXl0YEY1fdxZi9Le9+yYIrz8/M+cP5lrmpGIit0OCbIBiYTDQgpBTv++xT6
dZRxpcBK637DBKyvGbkl4DWJabrzyKdSERzO1a6qj5R9o8v5/xXahPZrPTUvnHVOzysY/+w/I7mg
CJhbD0BEEKAmM66aredaWmDAtN8a/sJuekgQZ6s6Jey34hPgbLtFbxdrulbZ8FZ7nfGKtnw6dpH1
sKPWW7LaTMprmF5Ke74W51dfe7/7RkZ7B2Ynhb3+N4cnIaZH5xuAG/ru44eb7Q5xBLQUaBtmdkI5
daKtkiV2lRewVE1S49vgebQNI41DEDzi1nmsVyjS+NTWF7i4lNmfkC37rUwgfKLP57WX3HCSqnbw
hfUGxz8ARgMeu4k/t8MuYx+4E7OcuyRvIh4T94kwwq59px1n5n/ahPJumH35L2svBhRZcUs7ul+8
gFM9StA1gp3t8hmSpozL/xNYMlQPZkBZ5VWiSF47lCc61UBz3qiGRQA2eze9t4z/U6aHTQbC7l6M
yfG8NDVwu3vLUvx8+lLmZS1PPf+IFfA0ag8WrfD+pbtmzXFlgYD+9hfM5j009bP5I1Lkk1LbtLHv
s1K5uvw/g6cNE5mrHqAuGHOLZKlAXuLzRpCJuHy86Wq5vkRiFrpAHnT/XmzO/9Whsm6H2DZ3780+
IrB83xVOy2uwEkDdE9rN2IxGKEGruTSFwAY5uIh3uSOboh0twnoxNvJcp76ewuWG7WhtdfS8MdBv
IIL7EYclkZITptO7bTom4IWx67/dN1UM6h+Kg/vciooTeTMUT4p9Y6sB2Wly7bDTpPBXGhtNV9mA
yp2hqginGZFJ4NcvFCyLHFQdJDyYcEE3QSXhi2HGWPqpbb5cemTwQ+rGQ0Ds13uQvAP0j1FiZqVH
SepapkfZlR0gbCkbH0INMhrArXDm9SmZe/T3XEgQIGaTpPIchZll35y4zSf1sO1Qjen1rwPJfrAP
rtdBlsks2FJzWJwax7VxtPFlCoAr/FAqw+tUvtpLg0bSeun1BDf2xTXQNK0UMuyl/wwgauAEb501
gTEEuMDmMJcxCNazMci0WaqGuLwDggnWCBTWb7S7JSHikk4xTK6l89XCqovVALdD+MEdO8EDTaxl
up+dNpaYuZklbixMsTrHhgnmJi5cHghvCBYhjni4gFi430KKjKbFkVwXdtN8EoiC79iDEBASNisg
6kGwX/EB56cB26uWk7EXSTR4AM38Hta3E4Djqa33oJYGwXUnbZig4ST5WP+6ewp/2EGMs1ARXrTK
Fl5xgNfAU7yJdETQ439Wgu2c9ImbNJj11T1oS5POnZlsbWtmTkYWWculY1BFVazJtnCuCjoNO69B
FiOS5FwRVORCFwGRHnOh4dmoIpTyE9I22VCECCrmsRlx0tEaEJWxQpnABbszUVfzceIqh+jQGeZA
pUMJpaTAEmgqGRrVW1HybVmLVLVqRtc/hPzQmLMhPHcJa8tgnpsnMRMRISmxzYfr5spIG5ADt6rj
PDZyzJvu7+Rf+VBj9KF9I9PDZlJpeDMEgDM9nA8fVDu/90mAZYCnFCnNvK+DRQwx8gO8MqLxyi+B
WSOS5hilfZ+Gqn8MFtyv4x1TQee5atPrPMAdpQxOqm/MkhH44BeQ3m1nSITzELwKz3cwM2HKHsHx
k75ST+SojnCUEG+MOpqRQDd7m5b7c5payGDvLdm2agPlbKOsAr47XcE9M/hT8q5vUvrgyiC9WSuQ
dk3HGyjCIf3OHBYlApPoh3LdH9drR/H6eTGF8kG9ern7wuF6jbEL7p1d5yXnqV+i871crezQk91r
liPXeXRDzNAGoBuLSL53flDhmPYhHD8t1m+Fx+NV+2BwghxdxuNTb90tObvNo8vjVp4Gt2u/znzS
3dQzn3Ohfott/lmQnO2orhDi1xjpCdpi6NoIwnn64/XNLS8BUcmWdvgnD16H42WHa42OidZuba83
hstc47Xs1o/yMFZR8VJgNcpMDh+eCerXos3ZzVDL/mpatqtuG4H6AKfpxLmESM0AorpBoq+j7XgE
DC9xG6/SBlXiWYPJDHqmOZa1tJR7rypCObYMgYVz93LwZ7ltf7Lf/tULCNC1CFbQHUFCoJwWj/v1
S4rRqRrLsiUvHvmshIlUE3YKyffRNq/ZQBXWHDAAhYn3OWutFJqTjeCDHr1XWu4ufLcrrMrVYcVE
MSzi5PU/QdLoleSENJ1m7tUn4ZQMCoBR9cUIDxrofFyDUlDym130XrohOs9LLy2NXTkemDrarWCA
msZ7VfRZscZzBWpCCu83DfacI+6WdwapyJpW3cjCnN1OjsvmBualOma5X2abAW6UyPTEUb7uv8gG
SzvSXVbxZX8ocOhd26LwzAejAat12EyFIrgGSsT8aQ/DMZsVsUEeTFMHTahcZcaovCc2f49gMWDS
Daw2aIgVCZk4ZLNRv194UYt1rt3IQ81U15U9b569we4jKXNhAof/aFYDm8gtfFG8/l+yTJZCLG8h
we/nHj6bZ45cgz9CezP/H8oSuFS5b/rDGDTDLqg/mhG9fNF0g3wChZFj5QpBsnCaQ+1i6nMxDOYj
F353+vKG9SfxtukV3pzhMRoh7OoPJgQHrZ522MubDkDV2Cay7lIQD0PmgmBdGmrliRQD/9+PmXfo
4GO7AgIX/DRUYU5RGHM2iMLkUfbTnR70bTUY3JcvcvcSYwVYfVVirw3AT5hrAvbD6e651WhOYR5M
qjdY2InHfT1TP9Y/E74A1laTyjp4opFHIjs/0w9SZBqQgW/X3MTLe6qxRj+CPDmOqofW4AzlfLsM
SezO/xpSmDhebA2u0y9LU/Fm8dHfj4E6zqJbSEqGpkepybfyWOdUjMnQNT+fW5urQcAj4Nd0gVRZ
SprTZ9zR7SlhjxNplVokhlMf/b0QYpIDMbL1gr/LtFb8NRVgGKyrmK171x4hZ3cgztUmJ+XeLvbu
kzy7qmGVaaQWYGXHYt0RcggrrbWPtp5nlw4WTF98VHZcEprlwA+NQhZnDr+aeToDR4sxk5NibQTT
OfbYpXlDj9xsivwoth5QfvOTvYiQ6iBhPpVfAKznRdgRzzCOGHhZTuYpsqSyiyF2xdm6lGAIyXxf
TUBKfZAXWXecN1XqmulOP2mYCXwOKxLkmNAL96Cox5tcxJ3MIyDQ+fBBia1QE2j4GF4pORiFG7rd
p9jue+MS14a8q657w/KLRQVA0EwqVwMXuaPM354xFyPHVWjxKRfSzvGkpXjc+MIEzIdw5FOErk4s
XwaccIz6c00pykOHrSSUL0eYIYUaQUJrFerFpoWp6fsLsQL7TkNtD5DTqCnqthr2/i7UKV55cpNh
6v4SBRH+ubY9f7Qz6ZHIaPWxAbsbkKLreOgfv1iMkWIVULnqNj4PBHZaG/wu8Efo3zizPOVKVnOZ
fnH+KC6kmkm50DdiuykeGYzKNaI3h9LbdOlYiJrxp6z5YZdHKmhhA+360KZJ3FEzqajaxmqaX3by
02gvWiyVccagQtq30kYH0ndIomEwJrsHiJONWlNE/HWHEikHkWUwR0XPcPTXEnBOQXiHUDsfuXoV
CkKGqMLEEYh3hMlrp6BO50OhNSovi/RZhez5JpXXaKHN/xJq/Rcdgex1BY1UMhwe5uLSCT1J+C62
PlO09uc+Uq9ZzhJBJLdiPN0hwEwwNPu6ML5spLtXK7Y+8xuvsCam7BgYcMj2xIfJKY81Bik0lrDh
0X0dbdNwEmizvHbAC4G6w5JGmsRZ71eIpPVIDpvDu21g8Q+wMvdlXlFwEujFLaT1kqBLTsrIWiCY
Fd8ihEC3A2B25FZ6ItKqDaqIW34tkGKhfU4wZ8PRSUq4oO+KpXBesbRbXSzgUuh9qL5LekQSirdw
RcT+vLeF6+0a6gRUWXUppFu/lhrECl1ODukZgIB82tcRlNTasT0/AlTeAO7fjIiql14WFyc9D6IX
+rDoMLQmTqnmmjCgK6mx5iNidX7oEvuKQDC4cnuHSW7c00LTVb4dS8H3I6Lk03MU/S4PLEB6uWHN
+mp5MNRjR6oEXvjL3W3gN3kXnbKhKNpqUvrXUJuLVlO3Zf9HU6F8zeqmbeesQH9AMkznON+4uxlc
UI+LoIKc5dwXEEqDa5aBi+ifVxjcYzKB0LlnajoJRw4eT5no+xkSr50Y7vMV4WFzgli9/96Ia+N/
TuD2wJhlpDztout2h3Psa7VH5B+oxNcUuBfpULLELBeRKde6qURHYfGNtiT+CgjQuYFxAfy57/Y8
a5GYrkLldntXd8lqKPxzr0R3cusR5LxW4HzlNGEi4EQl1ozcLBfn6ojXBIaNK7vvu33EZAXCqXXK
MPyn2ZqyB4m7EPYFx0xUpgT+Np/E7U6TnYx5m/EHIe5EEESLc20rOwvqhW/9KplVLBfnZDX0QH6w
pQ/Q+V6wky+nfcTfPVYu4hH0EI4dg5yQIoaoPA7+sAp2GI4dftz3dLnWEn73Z5HRIroeqGh0lYCI
KuJPPgjtZIAGmPhpyR8mJhuMzqX2RfDtQ2lAj11aGNMFC9cFQ6rQ+C418zRsNZAUeWtacTn/VTF2
N1GcID3W3KKS6yGRQW1mOFwIg26CPwVwrZqARw33wmSKFI86m3QfH836UUTEIspHmHkNiZg1WeSq
9cDzrD5uo3dCh1hAsJsw2ysHyvJt2p65g+mgsdd/R50BJeml6fJKNuJBerlR91H19O1Aqbdf8JdS
aV/8pzTXwc5MEwuCE4Vi1fyUHviski4IvsBSlgmC3R2ZDlVmE3Buk9m9AlsvGok+YQzfOD2CI26B
R/o03cy6uC0msbRt0Srm8xi3o1gzfz7wFGBjX10yc5BO8k8ptLUqmlOTagchBP4BL3QxYNBO8fys
RCklt+Wt0rklE3ZpGK5WppKtvU/5wXsjk0A6kPcBJeQVTDPWmKhwAyva5fJcG5WISBOigGLIIUjy
IxeGEmCIdKDy/cazOzk1IX86HK/2iwmMh4pZE3pLvc7jFmvyQcDPLFHgaw8KcNToJ4ZsmTF7RaD7
Iea8z5FtMdFBKzkmQik6z9mxciuasx/Wv2+TV8DFmszvc+1xShRRwYYIlxZhtg0/5f5XIYUe1AsQ
V3WgqQUpQxvh/wZWgJ3PPL79YpqRQqygBNKuE+OFNidZCT3RVcd8nVBa1ojZP9pTdLBS7EmrUtm9
rbXuH7l96bqY6Oc80SXK+sCaw/NXJzvIsnpgtSrYmGG5pzGpRN/SBh927x90TdXFWIuQ2Ed0C85q
C1SZCqKebzf7zUq9KgBLgW3rRRQvwKbqMdF2mysxVQi3g4gCUEkCITAyhXNhjtdidkYizSVQcxuL
j/H2I9jJmBwNE7vPNxEnnFHDVYlRxLM14CqaoUxANgSAKu1jUybPuB9RovWNQPWs2MstfzmxvAXM
ITXS9cM9ZPW/6EpgqwOb14kJ6G4kGMSeL7WDCrYyCSoeuDv5TWXvMGXqnT7FAX+s0U+pvqlJ7d8E
zbO5BWzsx7vjaz2Dq/Zy8Mfqf9OP/yxI050UO0suojUNbGomSa/VA10lcWfybMxttJFn2IOGEHC1
ZRDYzyJqxC80LB9f+t4JTNokzswlnCILw5ZdddsrIAqPaR/qxfNeU+vkpl9N4plRfiRYrRHXwHep
6JRD/qI+Rl5IRnv0gKgU9Id/JsNdGbxKvUZRqLr8qUlESRrE6nD/baSosmoU4T4aTyj9HLKFHTd9
FKu8BN06DKTvvktSw2zsX8mQ3mmpjbYMFp8FKjpUgmJ3A13XWxVv8TYE5YsxDhOcl5avBZCqiJmh
m7t/dqt0i+wuZknZd/tlgyViwr3rIlh4U/32i/oQ9sAltyyNIc3oYf0RpNG5QGhx1Ak2kyja9Op9
4kw3ORR4fM6/eMC7Rtl6MiD+Y+SCiS/59S9YN9/ewDUoLRCMfI0bKv+ilFS+3NJBHYxH+DqHDhQU
GEmqvfIZXYY7QFSNS47fH874B+mCBzmPoRnoHF0BA1jVIBAYuwdoM+VpRiGubZ+WYlU3Zy2d394I
GCdgtjDrmsW2AWe81dF/LE38+18B/K9kmOG0B16oNXafLmz/yqFDLwKvi9fwCYY6HZpZVv+9QhXz
V0HfgS9lhLd/G75ku+eePPzrLKPhk8zPQUMxdoUD6HEWDAGBXdBJForFVoB7ph9HlSdoPfG03jxM
QeNw7zKwn3SZ4cbTa3uib9gpfl5O/uZUs94X4iHUJGD2oD3+pYxQiixhr48/6gxoap1oV9JMcQZh
LUETRJ5w8HkqxuPUNh4HDM22THtNOawm3BagQt23PGusRLwAIszbsYzsiPTiMOpIsZIwbMLiBN/e
rTAJ5k9X/QQ54Do2aS7FrHjnt/SkGxrOabtbus2DaWbMBCIwZJZhvwPBAf4foMOJkNblTPV4RPXR
HUCSewN0iI2lKdT7VlpergsuXN8BJndrahKvglI2ia0bc//c0PPaJtbmTIY1EYZgFcOIv9imIyWM
fKNIWv2aT+oZp75pkh4LxIvFPLNeGB7bcAC+KD+3Z/9FGnHvkc6BeqF4zUKbQ4t4vYvWBQI1sfL+
FW04BX+aO6wAplcsjiHZ74M2M37UShS5B0AcX/TOuRo9frJC6FpgL8yr/yNrZGwnhpe7NQJzq6oz
8mbLidWtIAKFnvqMSJyvxu2zNRkkB51rz8Ji1tTN86bA9WuPLflNm9iob+AsMhub8XvaBO3/61Zp
ETOIUFtuHgMkysbyD0rkt5Cj2iZSC/Vxvd0/dnlzJFNvxbcPSW0H0n9/5FmLXHL3l+Q8QGBp2yzp
yxYzqBKQYeBp3bMbJSP4LhR8E/O6tXC7PpBfwYVZrjBxa5eIdDBYh3KL1RDX3//6xjCj09qFj2UW
kjDDjKRMlb6wVtlV8VvxxmSUGBdpPex/VbgEyzaD3GCFPRqIj9knf5jP4OEhZtZEI/6xE7OOu7bo
vWknClEhzU1SyrsOiWz65zG7TK7ACP94IOWJuFyWxkB2eGBzd7wtDUUKtYbui2dOaqOxuSeTAeky
bTwuhDREeGw2YCO2PbOpgXPtNwrvcJfoEyxFfZQQlbPP8bhqPoVjCvTbCI8Od5XrSKI24b+8VrRl
En4QILSqd0VRPb/FZ3p0rJfvkn0/54jbrSWRh/D28traRrpm2DcYGywzcbUoroPAWDDtWWkpPxU7
l5zx7CCv91+iBhZhwKp/1WbjUQoIIMNTN0GGIGZM0/UXN5NklhmAgbVQz3IYQeIWDe8ivmNO7heH
hK+MSK+YOurgKNLPOnxZOqXW6ypF7heghKnZQpJKXNjVhfqlfHmtfKD1yHpm1lFrR13+dzs/OVXN
d3NXByE2qwf1lK9hj13QAx3svffbPvKjHWkkskPQito7oNA/O4emSRkBLIz08F1r4Cn6w93rTcjV
JOuofHj7axvw+dpU21dm1ZY42hjqV0NpFg89EQqANMshRf30b1GN9q2+CciD16FKvmeh1syCDJSR
nArU8PQO1HccG4Hbz9/PqfdmdnUA8Bzyc7N3C1n7+nsPzeymKTXf6QZ1Acdn4VmUpA0T9surCCbH
MMJoDO02Yj8kOoprjNXpon+SVjdrH78ytWMF2ChuPUaiZlsYvDRoQLrq2E3YLV4qmzD4jVPZX2Eo
9KX60lrkTJ/laKoz3dLG/7CgVIxsnOqV8WPN6KmGvPYzHYFeLSuLvTRxVYAtahSFfmPJU/9Lx1ID
OHF5hcBnkH83xBlf6iRa8EQfmLhRbW60AyMtBx+iOyr71cU90iMAeoXIC/HQBeuvtHXTLZCmzjhG
bxU5Pop5towAdjv4fHBsDBB/L+Gc5/KRkr7mHpnDKRNVUnygoofDzLN5yEgHrBIClaerQFMr7vXf
0JSRw5Otj06xcLR56sOLZcdXvXcuTnfKjcLN40gh9mC+EVx6oRIVSIaH1P01bbBJQV3LgTH8/TjX
38y5B9AXBzXHxkCXaEFmvgCjDoCoRHB1KPBEW6EJjvesMVcgriaPqbWqiVSMJ2+KU5mdKNnH9THk
Db9qu5veR0T+BRvF3NWIt1zNE90FaHTt9jok8RXMyIb1vtPgBjTGcTsFuEKoewzZw2Hf2UMC4vQV
OnroN+Nbr6ViAnaWaTKDxihid4mYLojOhpDu3wT9j8pwRMNAdaZR0jbj2SShN4+CyefrnTg9gnYh
werc+wGjJYf+XU5RZl0IjOShFYixKLX5zKBGW9xYLyOsufGT3aKBFzClG78RxGbefGSwuCvclBKf
PTYqylRORoTCYLSy3tGtRpEkA03hPwtnWI3kgRl0jVHEjLR5BJJ67lsHrQuTyfsKd19zvuWfXdNl
jzj/XAxySlyriPVs9FlJ7sYbceEQY5T/dA1PrcnXytCgD3U9/S2wxPZszq2NpYjEdOU82GuCpGiw
0kzOJD1rkKFzgmJv+lQnG8dXE7C50PftOcXZTwqnsKLd8h8YtLjzfLU79NxLraZLTuOdBDiuHV6+
TH4lBtep4Fqn7gsCJ/hD7yvZhGsdxOX5sT0Y+zWukrkWXPBkjS+NNT6x/wL9KAU1udMc0N91PIrQ
2uu8G+1ISBNvf8w2Vb0Gtc+u/83iHypZKbboGID+X/3P2eB0x4f+m66EPXbFBqOgPGvLB1m9VEaF
MLsB/4KY8Tp96yLXvkTplJyAqz/8IIBHSbbvcX1xKAjW0hYNNMMppQ7cbhq8atmuqoGCWPRCPKyk
U6QbBA200CSBGkmLesms8X3nFn1mEpKzm7Sp6Bu7joaFdIOCCofFTKBcGklXKlWpwN8bQrs4PlVP
S7nm+c7hCkE3e0MSLcB4Yx7OPz9F7qD4ShvMgTafVTbKCbjNKhKuoCWW7H0WBSNK9taei2I3/qDa
7FxoaBV+ymeVF5ycMqXcfsp+uPSFJE6PFobWpnmm0tyOZY1N9QURWi5ILCxqDCL6Wi2mH5kkPowt
Y6fvu0l+177RnU4pQnKafuCJ7QsJ67ynQH9tu0mcjyianT6thJJm+8LrC5kl4sRsDfQeD+Z1NtJ1
NDKCFefc5mvaT+rV5NZ4oNyS6rFR0zVADcCi8o/NL/ydRyv2AHtaSzQ8yqV3uwhAwEtAQMQLqHCj
fdJ/6wlVYQdPbvDdUxhxQ8AJtBNcNA3V9gBjSiWrobEc+9LiTHFdKBk2e4EYDftwPoiBMIXBQzrf
V28BhTwUu1bP+aGIbVM/mlhxEbfeCuF25lkxvtvzzJV6COVmc2NPl2MF1TbzLv3e+/jwwdr+mkQG
15SA6Vel3Gsf5BpDDEAWmmjb0mP58n97K2qmBVMPpcqCBTaiSvKHpeL/n1j/hCrQ9YMurIook9dF
c1Mt83cqyV1ijitVOogGEUPkOxtdVaCpvgF2xSwpwFT7k9LCHjUnOIPaDDLnocsiEvE8uug7eMMC
74cZgyZgpvWkv7yvVIZr/5rIXc4K8tZmmPV3kHl21k1tamRkevtWDREvVZIAdOk3dgWHT/0Rv5VT
wwBay06vLP6lD3rZcImm03Ovxaut2ATnB5o7cTGJ3Vq4ae/eLsvFFYsb4B3FQKqqkQT6mWlO3z3H
wIywlUmv8Bj38GUAHX0iBG0+DKwjXx6dA2BBjid75im+7De9W4oJt89431tahoiFCTBVT2qxLL0Y
k4hSx6XiT/xHSvAaNp1bOjcDkyAkINY3w9rszPy0t1A231N4n2RrGmIjqTHPT8GiP5qass6CiktI
7VfdNWTktmBAKMueoPRDV633n3JIlwPvVRpLL+VZK8ABhoOzh6jS4aMYeAu0gBUEGl3RRZ8VXaQx
vRM0vnra7IXZ5G9eY+xzy0tCoAF2renVenahHmrMfUcX85AGWl0M35JUjxIKdvCat5GQVCQLf1bu
Fv3fE7bqALXn7V/BLRkitdmCatIThXDAW5dI+jeBBnhAgSqJB5idHxCiEIn433aAnzDawaEs4L1Q
9cz9Km89ylM/mbcA0KteZo+IuEdH+Ts6A9Cf6UBv1EyCcZKtLh40LNMnv5oKgyYA5wUXkTXZGeJU
Z2vTcxuflKsTQgul+l5bT8mfsDXwjYDw0mVW07I0MmiIIwtwk+QPeT71eJe1OBHR4OctSSEbBvCm
LTvyR0GoE7x4gRxFtIbYwKwfI+dCmYxwInlfkBuWu8368Oe2gq31qB3BwBCMlHAihhLZ/tLH1sTo
6e7ozRX8jL/oBS6u9U782Pur9H7DVBT7XbDlJeRn0WVKeF11CHnoVS/loCFMsu122RQxsZUPD4bt
vplbAi/n4K+l1tEhA4oM5knjgjbXwZgvYNChVvplh7et9tSbQO293cAQ8qncPl+IE8FWP9cyBwg/
VMd1CoVkbt9VuTQLUyJvnaIhx06Nr2+szFMuEvSvqaoXBddKqX/QtKIdeQKl9hVZdan9Dbe2ExwQ
bjOetwhzYHkNhh/fHESJ1TG4bOzwhI5tBI74g5uaGqBGwY/sV6OGaVPbO5LiM1ObuK1e0T2r9YIu
BGpFa47hc9YwXHB1jl+hGClj016C21PZSW1jRqk6ALoiJoo7BSQISwt2zZkeP1ABCSkvD+4R1ftG
wtSzq9JZfgnpcDTBLkQv+ffLXzGRQP6bAq4G8E6imaQK0yFaOfimd8uHPeOTxev2dJUg23t/RYKq
fyh+ZT0V1X8VzqymO1uEWGt9WyISJ92H+KW1WlhBwKd+097BLYcZ3O087f6Msj9wu1vyO2hg6D03
AX7bFGbcMxzfwe57q5aR0aOpmVX0HqUXnaODOdXD0F1jLCnChENmGJrBX67312fH8ZuFhFyBr/AW
jFNol9tcuUO1hFZ9WeZAPrA20sDm4z56urSKQgnQrhHCsTF1+Rj5cZHNvHOqT1fQWNjbLddzlC9W
saCEwq4DZ5VIMSWkaf8SiWWl7oER2mg2OekepWcZjkAKlo6xqbFV1Hsr4B7a+k16xgz3wc6sdTqy
s9xY4YI/mDUVmdYzMmGuRcburzF+uFlTMYCIqX4bbvgXnJN5VWkCmAyBRXpJugn3QUg2pyn2nkm8
iZFE3xqy+a3Vxc3i1zaeDVsjxvBGhuC7qTofKHesAT6i4BUbtN1eMCf5mWOt6759RllUV7p/NhQk
Q384rC1iGMNZIa9nY2VaydQ/rSB/jl02BxPnKs2GJJO21kScd9bP8e9Pzo3ShgWABP6AhztsFlPj
4SYVPJa+PzpDiooebr8TSDz3WscpeXcOhMxoICZzE4H6/weRGS8BVfst233WVDaOxCCyH2CgHRHN
lpOUShIbBprAsl2rLtTQre0pozzDvPGMqT0Fz1uwgzcVkLUEUgwUTeoBENyq+yjPjTXBjcr4B5mZ
UjVlTra0ljIqz1AQI3uGA8SJEpFOtkv6rvPu32AYwG5jJdI36w09J1VyazxmgewVcHjYMEsep7a2
ywCAaSv0IwogJEFXLXz0C4mSxvSYB7AsEHci3OFr5RgHHgaDzfePAgIBviexG1tIZdzfO2r+EcV1
HuFqeqvDflNUvdcsDlBkIyua25G/vE+dZeUuGJy4JuqWVb+Ktk7Q72zulyz0qAhpXxe8wQDysbdN
8UOcFzfl2IN9euK4o3pRu5VTM0t1uWZGil7tRk3cit4GUnflBbibwxaGe7hWMrPNwZmdzes6WWn9
bXMQx3DiFPx/uPopTITtxnkwqQUITrb4AH0+729AdvBDJzMu9D+/4bXWvLQ/+Silo2PyXa/KZuH+
KDBmbVIzhOLXkaVqfknhGtuIPJ5nKNmh3OiYluJMZeRyG8h1PF4VD4scDa64UAYCbXdnPI01VPt2
mHpYU8ralN0zN5i4XzgqlZJ9k906IiXqF/FxAQ77W6Tv9JfL7YZvLDdOdbXOV/WmC8k2XgITBnF3
LWy+mia/1tvSkJzhUjuEht6YiZAm/5bp9ZZtuAk4EncvK8oJ0Qej3/sPKZrPNvoNXJuerMRud30k
21Z1NQBv8KE4Wo34R87oYua1fkpeH0efjV4H1zQESew6pG0ZNArO39g/RUUYB7VdMtMmW6sBfEos
RKJvANlWzvnwlW75rEOPMbj7qjte0N/ZyHQ60wRM8It5FVs/bTDcPTBwLQUxT1LfNsaZj4CtVcu2
EBKroTMkKxRRnSDGwA1imDQNkVU0gHq+g6kSnjqCH9gpPNTB9KMchzDVJZ7ApysWPh+m6g05vp1h
MPEUcWKoIvBuMzSKWwiRKdgeTjwe30IbeUPv4K5vdwqbxAx8F3dWmgiJqJVAFp20YxVEmLkgkqm4
O+OKqH/Nii9GWDmESgKEQ9+0Ch4jDUPQf/ZbzlfTMKnbUIFXmyVHUuliw5ygusGaRE/hYScaXrR6
3KBr2qcIATYGqIgyowH/7f3+GuKIlXX4UW5oQA5lFk4rezUJTG0N3/ts8q2IJrhUdugJT3dBsFm6
k1CHYiGev/tJEyFGY+dRoimeCTK+rg4nZWALs7EKItudQ3zqyxeNPmmAs29TnFJ9AVgaK4jkKxgA
ofDj2FRzV65S5YDylqyT3MPwL84bjKlO0IRUBk1BinGrH0nZghUQpj1TZnjJUMcnMtFvD7HHX9n+
IaoWO0FbEnDpmm6aPizZcWp4+iRv8K0DYoaL8B3w8ovYzc2lskVeCXdQ29MEy7uBHmy5juqDvRYu
2Udayl0Ha4hOOz2tlS2DzcofkUeozyF5YjpjVK9Y16nMFgVlCidQtcZ+yucQMRBvviOS+PXtMAcw
dERLyqJmtDmquycr5AZrDGVvUBKvihgd3q6gVOiYBdQvLtOY3NhTFR3+8u2YkgPB/CKMID6oeRIh
njAQ7eDa4cAd+IEEvc86zxV+bDtrcPIZVA/jk8v2+5Dbu33YeGFde5SL2O1Erh/y12rFkSQdCjF2
+IgAGO8NbbXTWQE0qmVi8EimiVMOnUdxOg0cbjakdsvpxfNBomFXblwOc4rk5QsYLX5eBpN7qrNo
SO5c8esKA71ktdJtDbTzY/jp2uW8hcyEjI1Hm8SAEMKxOpng0BiCBUiwkzCO7TV6mjAO7KQW2Wp8
Mc6qP2JNp4qVjPfMD/QyH4WUeUYwqF/1jQbd5BS+oHD7Om+dniKcmYV1GtJiNk3M9gT/ziO6HME0
Kp3jryOZHimXnVqoNCsQrCWXudkzsQ7fVpVIfy32xNZxp6KIqog46T3D7H4TnFY0JOSjVTWDXfLJ
xTk/j2nLNRNsgQ9L8PWuNZ5D1aVtAOIYKbfN3GQjGBDfllRBdfDg8bMFY1uGlfQQK5pr3ues2+pL
8vNnOI/W5BGoA6OrB+E3g5Muyo1wfaWCAr2mdSZNoGB5+AdqugsndfPmR7m39XdKYat1REq7SJvW
j6jNwTBclF8C0RLr4Z7U0t+F4SU2gbKBp1Q6V19GM3k+7PTz+Kvg+plTN793HU4GM37rT902TAuD
/85pur33JCyNerhmIsS4S3orDcOWZjb6dLFlsec2qUc8Zw/soKvi2LVPsHmAzr3ri0XSfAYFq9na
6IUxHOSIZZ0vCPGQKYw1/5NSBLOeC/tB1wZeuZybnnn2WBlDAy6scl9t3T1wSFeTxf9S0Lx/CNq7
FaXO6HmGPY+Pp1lqexK+x67VCNiommY0HMBT5xFnSmCIZM4VmNSWZGVrLpbLwzr/tccI++t5R9mH
iXxTimx2REKeJTDP8J8YJTDbgCipLvFNMNYXJg8pvwUjjGg6N4GRNXoWOeBQkTbExGFZWFEXBpOi
dwYboN05r2fD3H1hvN5ZaluEJmITMMkW16sVXUcpv1jH5vdLIv/t8UIDodt5W2r5wkbCKmRkTT8m
GCW4RyOFcZpURi3VqG1H3gCppJHbZhyaeHOH0yc2kYmZP8oqwbYehUTAWBp4P1fcRb9Gw/rTc4zL
2Slftfc2p6PDF+e4SO5ikfZ1SWZqv64hQEbzai1+Fub8gaQx5xqjwj3jJgF3Zt3xmxnehQzcwSMV
VpMhlAyn1vypy1jq84fGvg3KqESMz2rzH98qvgFmvJ05YN4zN1NOMeybUutBLA1dKev6wscShlYG
Riv/zKOS1U0RxE8SAInUrm29gkfxhWhkQhmj10i5Eg1UUad7K49zZGqmXDz9K5JvBCUlY4dnw00+
KQIPbS28rfTs3KEFrsFXC9rc2/BbaS4PBmKMHtdSbcfaSgvG5+AZt7lFvP5LvUYgxx3rM0KN+N4X
8qq17hj58IQfi75/fToEvuOr02p6xL0moGbjTLo3CZhglpx5sf6UVNxb6Tfhin0+Va/tIxNNE9+b
c63FcI7HcyM5mdIMIKXd8KvUPud76y2+L+jjhLDJsNkEolaQzN/94IKrvhl2HssSv24XRiTClgLX
l8MjrVXnSMsqWYn1p7+KsrX1HDdhAcc3/C0wVYl26Z7LTGT1oEG7oEvE4St+QkoXU8M0Ph7IG3Xl
GsikdbHSz+sjUGMmFewTgQS4NqunL4tc2MK6ndKXAIc0pkVcxXsn7wjH+h0adbE2V5h74QjJQ+8F
H59FHaoo3Rw8qdgHTrao0bmdgJbCqmBWRPiC+MY9ISW0Dn2RHG97HoLuNWMeLZz2yJg1+LrTH9pE
iHPFC0V+QrOOkabqFzp3Olnznw13ysuCJZxoAbQ9DBz2lyhnAx8AU4A+w4JHiFvOHwO0yIfaQwpP
8Vy8vUH7BoxIGqbYNk6ob4wnBfKvDeXksFH++3510HwmRkohOPdDfA8MXxWLD5vp4my1RpDm2nRs
dt0iJRhvUFhrqqBphMCFX0g8n5zmSda/gUyFGir4aP5k4FvE9gVaX7ByrC84/n5Qclf5UC/qy0fe
NfRpubmVMm9PJH58FxKMFdVmdcP4LX/lEoRYU5WRC0+88ivGHkcQAVIGnk5+XBlsfq0YpB3jOoTM
3K0AOWgFUGtIldHAWC6AZtybNKukxEyzo+wzEGj5/yLVypSwKrkxXKlAQeqMQBKxkcjIODT1s+vP
PGdRJvV5rXxtB9bSjxldQT6w/K7ZZxFS7BfLXXm5QyOg/D+cnb7X198S57v2m8V60rEElbozAGeh
/JJZVGXCl40v57+9839bcvkkZH3jOD/d3HLRwrhWPWmsNhY4jNq6KwYqJznT7JiJ7auUDx1MRfUB
jVfjdUjvMsO38wPvh6HX0OzI4w8jhKA/lNrufKbhjdlbCglbovzwIClyLAaDOEjm12r6PMtwbHmS
oRjGszCXzspsOI1lJBnd6ylhuu9mEjERTtBd3+mLzvOae+2k9VUKDdoxdrh07jAYhDCYrqraQUWP
DlOiJp13mUwJHYJZX3V9BsCDTVvcALUPRX6J+KyUjJm9pUCUGr5bHpieJjQ+hhfLdsXPlbCeAREV
WyFi8yuUdo/kjq2Hrq3QQdsbFwzn1jX8TBu6oTHX8dUS7x4/Qy1QRKnVm/4J9else5LpHTd7miAu
0vvKSm+/c32JPyYLAYx/GI8zqaDvZvWmT9y5YQxUIduQvbcNBPXJMcuh6SaddiEqLbSYLbOIouNR
IHvVQuB0+GzryIbi0slbj8zfaoUP0e1PyBhRU83bKvpCyCr+4TWPuU/2wJ/hlSXHw03Bp+zq7hih
gdXLUegghVHfeNWXrc2oMLNaDE1MkIUKrr8XWRG1iXF4X3Ht01Jv4TDcXOm/baZaG9MyqUQEUDhk
DGi5xb6vCbWP/4Db83mABE3p6TNYskb2g1qvdgkq/t7uaKoAt9zTafLzm3ZIvVr03dSBUWh71FUp
OdA9YtNOPv9j+Sa8WI9lUARVanXZ1cAxPHyWRcfcXHJdhcev9S2Yf9N7u1Ge6nB4EPXcNuDFFp/s
mV8tv/+eXOj/vBpevC+oN0RNTNFofFh9utVnKzp5dNpgd/bB7J9DwSDDrtTzTygrbygVOcj/jS+3
YMcw3pN9jJHu1gtw9NdD6ZLOrycAKtQsElwO4lx5+Eul0VvoeGSS2jDptjEDJAb7yLVE7Os9P8zt
x2PLUP1s4RL6buljkpNT7pYYmLUABtxsFVY8ZrMZtUMJnL54QglhJOOCk/gpYiBtGYrYSV1A/Nsc
6UCTAcLOkEL8gg/8B7dsM/HQavPfC0hZ7koT7EjuwjWnUmepZ7xDW+L7TJawna0x/AeSA3VaQgAH
izNDPZbaQo6K3piEPVGAVeNtFn4Vw9RCDC5Q19fKod44AbyFSdt8cBhasAqkh31Mal8ZaRYXoCRI
h5xV9zrVn7V14Q8xMLZmDJQ6TXh/MJeIZYL3VM4bFZtOQo8mLoPnaOmpWRxxdS89JnJ9tY75E4HS
zouKYvaUc1N4VW6bigySuCkB+MsHAgSxkpC5rpPJkmqH6+PdoEODT69YBD76SVy8etnq45RDDwdd
29zufzZPuqugfpFGS10XKbimNqN64Hq0G0YTsCbfnJAMbp+xC5JbL1N7De2VjToEM31uesfCEAY9
qDvmLEW9MVKpz2gTtcW/5xHi+XlTkA3l3khCMXIJFbhw1+Ucx/d2rT4ywBTHPTEB58sx5TdvmHr3
nmkrMu6Kr4TdrZfa5jHssOQKtt1GVpW2CvJpLr4Y6iMP9DUZxkb0aai5H15cQcCVySiGJx77E66J
Uevw4ZkJrlqtrEHX/7PctU8O723axFnDidFpd0yQnrjTHtzboiFnmPQ3ZQiEA9WAVcwNXBIXT1/a
aSu6Fs7BvCR7FLqDCBU82JwJ1Wnuflxt+ufz7VCenkNrszYGWJynLrWEAXJ2igM3ZCVpBQ3e29x6
vQ5NKConEw1SZifBC03z2SIoJnQeJKPqEo3reME4lRG4ID9mku7JfUSKeLlfeRr2wCozPYhcpcoy
YpOq63oMtTBuR8PPT6/qXJddVzGiF0rJSGinHziBzH4kgj3XGETVGnu3kYpJdNMd9bGCcUeW1MSa
BFklV4uCnUPatGRWsI5I6v7dqvz6yhUHGa0bEXWBoLKk1Ptz4xMDovSYHIOHnXtwRNRgX/+IAHGI
W3q1J3RjvKNPI/sqA5FsaLprWZYLNpUHeQubY3Ptp+Oa/TSYMAfzSTAjqBp9s/Sp16C2wis/O9Ot
tQcxcAds2+0N8lp4Y8H+2ZMbVsiXX/u8CV9kluJwIFkx9BprhcHskdb6sHGeJo/f5bUPGCBnyrh9
/4TS4lK2DtaHOQXgK8/DHxusGTqAvxtQs+jY36N/PO8bZOkQqQ1g9PdRvwJXl7Mxm2sKoosKH5uT
bGVjmytfVSCNd6OlTfC/Y583R2pHGp8i/75dTRycm7WN4gUTHGRny1eg6dOS1PHbZWiPWC9Kye+j
tK48eryyGDeN1W4Ac3DfeBTIC5aDmLiNdDYUVe1C7iyeRvUSpY0nH9Bb+XLTWQh1RZds2yrTe22n
VRIS745ZlCYf6uCrRkFI8KuWeADG+//HKVfiDPKe5MSSNRCXw3XCHHVVJNqAXN7HIRmwFE8XrQu8
Op5ysZ+/DzpzlUZmgxO2D/T4M3E/Ku4DVqOkp1WSDW+0LHX2dU8KmQApvFpoNK8nyaipqBkC33dT
uigwGneAu7WNTSDORSXBvKtdUDWeNbKIhZ3/05L5ByVmkPi42oTCXkWHu3R3gmhSmlLxOTZoC/Rv
khCkJL11tqgVhY2Clz9FGk1WZ8p4H+JKKow+JL6y8jtrTKgd9fTpF81WvdFPVW/s8CSpNLHTd/54
gB8w083Sf3V0jxmt19wHkw6RJA1fUMkbFKN2pYF2rvxSkdGz0U6kd0nsRA+6bdkcAno/n4Zg8SEV
RwL/qJHdpsSL5lwmeEgYDk2Rh0turwy3YBUn1fL3duCsl9dmeDls5sBAuSS82pI7fejl0wCctB6P
kvUicgrYZuoWuk7xEz+xi5oNgtTQzGl9tmBFKJCoY/E6R//xR12ysNqLloSWA6HUnWo4p/RC2nPS
6T35fzWbQxHGlIWHz8l+XN68pg6oH7ToWhe0BjHhNyVgwEwx8NT8zoIczzhvf8hF77tHzcN3ck1D
rGkKEszRClOmN+h/ZE98BEd7r49PT8OsK4OA4qxMxVEfIB/QoKObWDYyJR//JiP1AR8R0WXfL9cA
Cv2/DgvYJnGhNwWW4T265tcQ8R9H195yJgVVDjJgPL+1gGJXSN0JB4ny/WhCqabwTcQ+JKr0olwy
Eri0O3Av2/y2JVD6sRIgm8otlQrM+Ht07Mh/oKo7Vnyi5xFWkI0/wT4dewAcImYJ9Ec9YZiiQi5F
Wz3YZ2yhFxRM0T9BESSOwvm7NY0sdY3H1GvmggmRcfTl1QR5eE1cEj7gQnR52rW+FPgkhvaHaOTK
99CdedJk2kryTpKg08gyvg3NMnizHymXULXknOftT+Mcy8W5LwElvS0P8yDImUH2JMiVHxaYxwLC
djMMzKSOU/T8nzacs8dr6EA8dnQkIrMgumZRYFIcKDcOuaqv/YYiFrPyUs1tEp/xEdalqfs0T3kA
ad46FnFlJsGwwVe7Wj5KJBkSnn2pVB3fyMK2AvpZSm7+twYQcVRCYbN2J6hFVpvB0OWGdHj2YXDm
RnPYvGEV0MIbETYWNdpKxYMQZETtUIJGMNrmRRZG201Q9eBdxf7dl+FWDzKPvaTVGLWwI+eYlraw
5eLls+0ECP1BKASzQ99Ljs7TShfKeqabZq0bdl/zI33LPscdEPuPYyEaEtdwYPwNCzHnTMKws9hI
gd6UOWENhxTBItw3vp3vqaItTYnVs8A3bVD3J/7n9/Q0gjnxCUoYHG3luuqP3QjViCBUwHwFz8S6
QH9m4cpWWm4coVcEMS0Nf7tyZqziM/RZhzpUnDqTDUaoV57W14Jklr0K22aUitUhdDoGiToiNjNr
ntMpFh6dS9ESvSj2r02bQlGffa4F1MmlFDTvsyoYSaQi/SQ/7M7AHgz+K/5kHnyiXcUReFMRGrv/
5IbNc+Ruz7nYq3Ev4OnQc8mxVTu0Qx/UjE1Srjp2fVam6UkvpYa8OKGqy7nhCeadY/29hCzBxy+x
O2y/+EfcdS0P3IUdUa5ezdb8CONob8x0I5RCNuXYCHJJph5tpmpvNgnXBm/8/MJijPLQws7kl4Cy
FL2oNJ9XyJF5qtgbOIPaB0rjDSDB5hYIUrrMWt+UYTzTSnVVuDHFjQR7enbvSeG74t3khs7lmaol
mRTvH2ygXSGele4jMeLuBisGOe+iip+dnEHbv1NuPfTKiQHVYJdu+saKEc4+hg+o/ooVrPwO0jU3
BriEgpmCcVtfp+e5eRhsRAMI/W6hGkKCA+HROPkG4wH0ys8dwrhIUqnrjxSqrtoe4elf12OKK8Bn
VnXm3zRMpN9wBhATqvknoC9HhCzAUvsq9yPkMsoaeBklwDvvIaC4Uxud8sf+mG1+kCXBadptHvjy
6U/MAGRELIK8CA2oX4J4i/6pSZKDokBQvQ3XyaAC11m1sAUD0YQiHUXlZUBOCVQE1E7Rh6RfoLa6
Fd0H6iFHRVPhGYBkDt2jrWKsuav5ndd3KSvJr9g7miaDmr8qXnJEhlDawdqjrwKjVxxe0uPn3nYx
AamAOqR3t08c+kzbF4YR/NoxpX3DKNMsSl5RpY+RM8l6g/fDAI47dGvPTcJs+QFxWJpb7MJhkqX0
bSU9Xi1fTkWwL3aPbpOKJ1yhPstRuwXlvUbRoypOraohUe0JDtDf1QT/7ChBruQXdGj1nnJjco+L
iM1hnbU5dkkxLqOHj76VpREckKVplWW7wjih5jcOuD47Y/PCx42LqkfQZo2vm00/yHsxswg7ldfX
+MhrLJk37FfMYZCUSmpAymOevMruRDd5kBT/Ut5U6z51XqeizUQY4le5EgidajGcr+n3eWy1uAOy
kAyLpCjqflA3N7S2/EXLwflUyam51WQU/xs8llIQjsBeaiCfP/m7UjixVpa1rTD/YWKbJegv5xNN
V60LPw/tsnsXmIGUC2Kj1cbvaDUHoZnyG3NUniJzhclzRSrD6WScNVJOZijBw1x7DUUaicPFWvzq
PxpmW9UmpMqHX1eyuIKPv6m/hB4tP2dQn6kvztwJZN5DZCDxIuOxxXVABdOGUf+krqnnNX+ue87m
GzYxwr46W86xoTuTjT44I3NndYJ7/AyCC6NpcBXomB4C+pExY92JTGNwCAEpfHUKZjH9G+70Qngw
T67y0qeoZ1hr/j5nSURVogaIFVUmI/+ow9tDMS9rVsUIqfdn/zyfmW4ULwtHW/rHugLFEmyzV7wL
kecxzT29tCnthYAqximXcq78kGCBxNdxzpuhj5z+/GlGx6ulgaL8Av6GV4KRQpX+/LTvtNuuQwHX
Kz30xppCFMesYBZ9bYNh98pL5MsOY4CigwcMqx1wWBMUteZSF2kVHvHbEMIN7M6G7aiYfsYgzYAf
h+kkoltjlypjuMadoZzQPnWGlFWV8kbgwBlJbsoFB256ursZBGktG/S6g/DiyImTvo7CqiRE983S
TV7SwqZWDGIuAqDMzNCVqbuojvDDAVvXwAmjQBcSbgJxEUKRnDSuqXbCk9Q4p1OmZBXQyoAwuba9
ykKseyH//hoOsjEtyVjXpqNEH2SDfqbMp/rOMMLyzwdc5gP5PvbssePZbqCYRQlf3pAs9EvyrEen
Vub70a/WMhgQVe/o8JMPWXyuX+rJOqXgEe2RJ6Pcx7j1IpMYqa+h3G9isvxW8/H/JjrWkhMbbceG
qrSBKpjec5eYTSmVP/MeDxlxmye3ykGIPe5UZLo5JUjcRTtQRGufeU27mWEvTW2mHXAlJYgSOwjA
x0d9w8KINaBDfwFUnVwYM5FjQH1ExlCZzf+Mg4MUNbRaV0eS9ZlJLDQz2NK6AYM/MwWMRNIpNzrN
UhW2E5pp5CaFWHXfSShS7uBF2Bdx/aD8NlU7QOrYFPMbHsBX9CQ0SQp+iMUwRZq/Nv6QPr32raCq
z/IhFnpITBoZln1I/pwEIcpReb8KnaBGmXIsgu3jXUzDWntsbmaGwvMCGTW/9Lt4eSxfBsBZGo3m
el9YeUdCDa2NQSt9nwP+DBB9K46mB2SPKMvFQ+HTFKksj7fN2QbVKkwcvqYLjLIXm6vWXv3z738x
/ckrKmIn/z9SJP+/EwnFeQpocqEUY6BqmkaXp/WKhTMsTMkNgGEKGaatggilJ1ROlCQLlKO36CM2
lZNyLf6a5vwBRXYc7NkARkyVoI/GF1cFClrjyKwyBcUxojkngHiisy7eyWLGczgG6XEMjh1KqExK
VFLLWeEp9FRIZl8A0svIwn+KLgUYTVsypsybNIs/dUk9HtHr1McJoryQuyrXO8eIrAmbe4warITo
d9ynD4syzuAhZvRb8ufR20xyZTn1kPTC35CqenDj2QEemsCRSbMhfBPAxewT3YgvIsg7j5bBMSv9
HwSNiB7yFYe/2p3Cr2MQZTXelvsWqsrlTFIkLHwRyxOk3Lse4u2+1Ks0RTE4SSGzIRHYjWPWKCd4
kJ9P14xa8gKCgEfE7zuPPytNb8MUNpAdyewh9YArAFl58JHrRE2HvGazfUNsHjER1tWMAsIQ7b9E
tEgi1m8pop404oFbGLkGhe+Ih0O1PUDBZ7tQje71wGSt8GjLb7jSalIRFWmIbmgJrAhLMB0rrneC
somh2RZVWxd0qscIHMlhY/bhbxIfRIRS9UHzRKH2ccmVSPWvXB9ZQQomPZqSFNCqvvm9DgrO/2my
d0IqV4ZT+31jhzB94J1LatCNDOk1V8a8cidnulcb2V4MzFR8jUbKrwSx51QhmdaaPvv/IfcteK/A
MEz0D6hOmfuYblDDJZ8y1SMrSYPwWiapVZYx53/GyyAXpMDod9oeaJwlebLUP464I/yT3dN44tgS
bGV8U19aVPy+KY6Nm+BdqQkfu9uIe6M4SGuL5f/nzykYStw1DYVoBgpuiY55nIc1znIA0pE5EQLv
HEzlm3jE6o6Ar4ccIkB1pAPkJYxkeRItfxpftooTNa5/j0q1atm7Rmas445tzdu70/h6k6o54dp/
mo9XDS7tpglzqE9+CNHR5MICtnAqiYiA9IvCPiZIBrSrvhqSM6W62Ao3ncdbmX9ndt47qvywqaPD
VWbaQmV291tvGP30OuT5ZEK4XIcnObRftr5D5cP4/G2T4tCgtis+4lcnLsVc4xBcjmhiUSB7VLs4
ACLG9jsz1cmgJ93+gIPa5+UBigTZzcy9hCKd5ARoC/xpYa99BYBMtwul7R4JvmOh4O7+QJO7U9xj
kVqj/1TQ8bZ32omcToZdgWqfhXd+auZqYIeEK0X7GqSJy5QFrfIEIcKDT+EC3eF7uVyJCxX8E/kv
RLTwCxgX9EVGGiXy0zVfZahrfSY+szezmsijxSI2x13IEwjnKU7mPM2o0DsvOIN/yUBND/YeP5kn
DRKlwFX5Rum+M3EdxMCNyIQ4pJPTMFW6B5XzEdgKBdZuovlFKj0D5aM/cpU1auRf2bvo7XZP5vZh
2lyzeepMI8YcEMEsJgUuGJbprmi3GgW8t+3BGefI1Acz58pl4BK2Nn1vbIZq84V6PdLEUNNNJen+
tgxAeZImn6mDc/vAvYYOrmXPoac61q79hDmgSAf4/Lx1KF5Hbpg1KUKiJFbg+5/nvnobkLLlxHM3
lYpvq+0gY6nGlESCT5t4p69F+rlzmOmonwbhfxMEYGaKCq66usZpzKT/OACkMLJPTeJns9NjNeak
P9/QQChUt3KUFmFYGxItnDtDkJLGDb89UdpQhUg/xCgyXW5Bu1OsOgDY22Vlim+p0A8S4CnNYDvJ
D/wcVO+mxI38hAMUst0+F8NV3yYBUR2RgAeyYDxZODDCd3h+veUJVqDSnQGTvL/PDmdl6hLjSngc
HT5Sh/fUS8V1/MvrIVHd86jprKNKjznuZD4Xqx42W/A6YAJ2GP5vBZpMANUdG27KlJpNYkSxH3hM
o9sr16GVfmhPOdrXqr2CE/WUE6iOWXGP8FegNa1oxUPocSG/Q/kcTP7Q6ZseS8WnEzKXYZyEKVvr
38DCAlryxM+TNZCQo8RAjYN8VfXlKzDPq/VW4KrVUZi/bRZeAoM2hzHsWx9k+MTOcmFALf6nW/LZ
gPKzloh4/L3+5BCNjhkKILmWRM84rYCrUsnypgmI1xgED/w/RJtanNLlq+1ucwej9qPK4thxia6K
2tMAtBkALPbRQd6sl5wJ/CzwqQLNUDThgPy8g1uHXQTkHnoY1uWP93RWggDbLPka/CIAWUp7buTi
WtOmWGS/lLewZLzt/qZEB/AN4yFkHeONaX8MuYD4gjJlzYxKD4t7xM6gH8z3sb8QPkce0NbbHmOj
VNKA9Z1s+F6SlCthGiuVhKqCPj76e1mq4XKlOOQYoqxvOeDl1nbondpstkz47S8HiZKJy9iDInfP
d5+bIaXf7b08chaA0eDR7YCHvfOm3P24ED+nTFb+1JPuCsjyC32HwSHGahp2k5XIA+Y3fptw8k22
KmRF4pv4ECutpp9fLMFjk/kQg1baC81hTwSq3nwwFNtg6kvvUYLffzc7Mtnm3xeIM1D+i+ZX5Uyz
ozbHk3AIgJpnw4c5wYP81w/pF1G+EYsPAYtU8x4NgUSQQkpiG3h1obV0tlK9cFfHQR9qLZaFIUy2
zpfCb90vZhuUIspNNcOyjqSa40+g5FNsBeSWLGxuXp18Od9a77qrdWQRhsI6kcKFQrWV93A1s/bY
+PQB/DFhmghcHXl72F136vCgbdxoBPIp7o5BHrr6F+ljn4dcXLH3MU+8FKgUwFD9hbxHlAajZOZv
BBy28vll8bmQDYS0FYpXUXx3EU8rWzFgd9sgO+OfMHvpWGMDTJMUHcr8NDjO73SKdf/YYJCecYJw
h1ThQvmcx0UJJ31ZzsXpK3O1ZEmBFgeQNE8svwTyUPLQ1zHMTLlJuEtwv4sC0dGaq1eX3TTcSXoT
wVU395R60YrtlMIA25VCMTGRdbkj3zg/h4XJFIGoZQginmM982zDYjrqDTNswC/C3KGVAY7uSeez
xZIEQiBteRpd+9UMmABZD4j3KG3Ocvqn/sSnpjAg/Ma1NBRyEcHXmNgCGolGGSF+hf+/2D5L6g5V
omDDia4SGPe99sM5PMz0UW+DfutO7JT4q7ket71QwTGsQf4zDR9tTWK/MEnF33ABVgBDFcoegnXZ
d6NllrCN1VJ6MMOlyxzXlfRoRPqpreKbpYrFM1w6B627+dfwmqEt9plwDKXeY99rlNs4jGhxyHaN
PZS3QA8LmocqRdTS0I2xWRq//XK3Dgqt4lNG+XDAaHwbkmBaZyaZncMRk6d6F4u/oBARDIJHzOnp
iLkJsMK6UF1OS10Z4nMEP9Dkdytp893jvtDPiWS25is9AMWjbfxi0M8uHaWDNfYaBTyBHrKMCXRR
9uY0TvhyNiwGwBc5h0SmXcxFynWGHoQl8nhXvThRSsvdcIUSHxKHvuJLx7Xz6AB9/9s2Txqr6ZjF
PUaKo1OYMGmoVidD4PBrwsRUXo5bRlC0nYlJyWdoC2xHzDsw0QVwN1/Kj/nkI0zCePIX3qAiMy6x
SvV4Lb/Wtac00WgP29I1O4ODG02STAagnKDeq8yDCMDpl050oDG9kNrUfpLTKN2k4EDkybUvx7il
v8tg2k6wMPkRxL53YYmmBKzQYPk90vY1A5mg3VQSXdsb5TKHE7uM2vwsYX6A2uBSBa5oOAWglQAU
hF+sECaI/Uo1+5z0zwF9zPYZyca5fOxpCx6VifL8Ld1kBEUyS+rGJOPeMRPlkYrrTgUI3y4M2I7E
810VDDT5p4ePae7ArWNm3IQ2INoUHcLShL0FnOAGvQXofwhw/ffpnIWk25OTrrj7iuY2YphQEKZg
z8H0lBVO2756iaUkHWTdhggMcuzjnnbJ3vX3zV3hzThF8HuhUcI44yMV+3CgoJek4Kr/PRUlsY5X
3kuwjfm715Va5KiMt9fM2Is9S3v782Cit3tW/P8CxFN+pSIkozzpyOeuf/KVxD2UHJDrt0i5OWW2
lgo9tBAdGVbvqmrPakTCSt9FsUzuXMa9RtnZ3vzBMmxrBoJhZh34rAlwv6S7Zr1el5UhiDrpiJKw
O8dy7rPN3pcRWgBHMQBhGIYJMOvCgocm7HFDEmQA7fvmc89EntVkpLmWRdrSRIsVDsrf2jKk9qtq
1I3cRFoRujMrF7J2Bv8J+5rJ5TRDtwuDoregLCXVUQtDlKRaXT8OO9GHfLZk95BEhDNw80i8xr5K
2ABQldksAaoiTvwT7lDi7fmNEWA+KToD9d3X8hk+Tmvj2NgjbiaFv3/X+ASty0JMHMNwLsN5vVzy
lMusK7U3o/WF9OwL9LJ5a1iTsjeZ2BwOhZOXNQxyARMAqI7rxBv9uYjpgzgOtJyAW12X/VkfrrS8
Jisgp3sR20pISMrOvFYNS8X5Yr0KTKFIBnBzvH7NLdz88QdqwVm4jOc7//jiMRsekWhvKBJiR1Do
EEd1QoB1qg5peBpWI2cSPyWerLXdjRSZdUXX6qCc9QIr8Or5ScIjueBATn/KkVIrCnMbmwCngy3z
lW41ZRBTObT51/PM7VXbHgLPTrZKnUYMWbnLrKFArIO7sMUW+MF2S4IDFJJN4NWKpR3Olf+Xvail
adlbNEXrzzpkBjjtSu7uz0IMc0ZtDWhEb6wcD/fk+ED2hBM4iAR2y4rn8uHBsdgP2amZ51F6AtPr
+lVkRP6VdhUVk1A0JEAL5nWk9ST5vM3Zmz6R737IgzlgtQpTNrD2DUhQRHe4RG2TbNJ0vUfoFuOz
WuDfKEjGw7FMcida/dQ0T0Hq6D7Tgh2eo1xbS7TnxF30I1JPTXstxcfbaw9NqdIJc97IEmpp7+21
acaiYjD7hjYqD9U/TdOpxCvdtVwahKFS+eLeM3Uwx8qaLkmPdAHbDBqcAvy3KcE+TBssbmZh3Cpp
1qmFPK19xKmy8+56Rh/mL+RgEav/LKWHXhiVf/EF5KRhsHHbWFjcP6UI8ec2+2aZV55XqNmDyJcY
44wBlqvsG4FjmcKHogOlqetAxJDsC3jeFtPUdMQTJmHNKIxYdWmqG1lXDfL0G9wMJevnjTWWkLL9
D3DkjIxnOKKc96QE2lyC2YLDnJqHr6EAWkK93mDOj4k8BXE/tsSeq9S7ioWMIw6fwqhacBSScQAo
J5Gu8XxUDMT4e6N6Ce2RS5vscJxYHfAm+qKf3KsCdKVwdm6WXyIXmMCVXqJcCQI+uNG8YwfmXBcK
N5p7UMo34DBCGJ8dhN4+LtpBPIVP6J/7rkQCqnoDM1D2cVcEeDToRNH5TSaPM4lPuuYtbNKhH+YQ
BEjdWI+FBJ+ARRE268Ac+hx694BPPFz2WXbd6p56PwC9W+lRBNg5NXkuh4QgQMU/GQZZhxhFwJIm
0rcYGh5K9sUNJT/vySPPyc0Me+b+Y7XZDIt5/y5jG2UZnMvgnUzCOQHwJ/NzEwwv33S2+gYcxRqZ
eBSf3ON7tf81kxsDl2zZk2M3MjYxmX4fxBDozMbIOmSwU5j2JdracAvL1mEBVTgmvCN7ixZ5MyTT
83EEOkQdc1gbUjZeMTtzuKq5Ctf6+YhfrIpy+/qGMokEQ/VszrqVmlMy2PwKPiwpyeS4Gar/jw71
90UqM9tc3z4iMLpmsPg+dw/+5tU+Vutb8wQrzZ9HskJxQ1RgB4xdCYboLTUj2p2R3QWELvEZxvc+
LpEVsjU0LtZW+EmuuFfcEd+WRilmRoriPkE7EXs6HB4VSk/UOWoFK43Jw1EHfrrO9EHtWGQ+1UWs
JavO9kZnuF9kek4J5sDH5//ZUNXS0OL5A2Hg6Vf5nYEoOoBfrJpaHcVNUI7BT1sIBFsj1xyVZvlJ
FbhYCt7af01Nhp0X6wXFL00Q9rnkdFVYXLxdzi8bm6PRvi8JLFjGzG4Y5s1ePXQbND6CQwDUPq+n
2g1CKfBw4zNk6PbpA1vIJyA5WOeQzrKXNP7nTYKfGQa7WTwznipE8MkpmGxoD5hEVu8aA/RwIShE
0pmdvgknotPuKacM9eoqBde0KY2ITq+DrBuH6+kcl6pDNrS50/7LE0TnK50XQV0Pda0ZaRInEvRN
LlmVmb0t9f7oSyBm3Ss6EbfYbF61EzXotEHzdbICKC1VFHm1K4eONksie/LE8mTym1V3BcA1z29a
Q10Jd2Jte0EBS2tROKqOH/JhGY+r4jS2H3tvdMIrC67wQqlPvihAn/98u6rGVAUCrhu5NEV/fIOg
sGD3Syfcw4nYncZolcKcHu5hEBkV2NXr+9B/dfDcFQMyZ1eaBMbm4M2VCg4/gNXnbUghhLcPpcO9
B/qpG7Re7jP6434kGLv2CeJB08/7QznmZbeY36S5O6JIpGE9K4THdRJ5tGBiPMyR8QgMTcchKKaT
VsMtIlJldRxjrh59rQ3VH+keQU9bLlmMfqY0A1uWRSuD50glm/NeuA9NwVKXXqaqQoabXNgZT60v
oMQkYwxy9BGFCNumaSp8XkPIFwypPht+j6a638v9dyWt48OQEeYwq4/YO5KpRYIvLSDCci/ST3Eg
ccN5pt0py6UhYCdvJiuIyBbgQ3d+hGq6Cwf4Yc2Hkm+WzJQ9N8HfYGnCF82Plx1Jrcm07TNDzMLj
vCPQF+GqrDu/FOHS1Iy5O7hC6xFf9/UK+zr96Ml9GiJlTQrV4/GFZE4qgwVKJcSnF/V3jtyoODDU
VcNc+RfOh7rw8pFfBZf4LVeByIyLVttY0xI+k1Gj1XBPW5JOW6Ihp9tBIf5cNxceby/5R45MAS1j
+L9mCSk5x3jQHVCmzs1xSXzceCV9SiA3WtAUSpTFNKJPqNiB6G4wNojifF2QI6KE2K/HajSXF12T
LtiRQu9co1qJUVw/f3flMSfwCpJa4o6iMZawQTE0B47mjVy6QwMP/uUJIi/T2Zy6NTzKni2TeUrm
WpAmWu2MHJkiwMHCkab9LMnbcvQJsMW5HZ65/4jrHuQtJHJXuljec8C+OqV3QC+puc0V7xdohBOJ
cxgyNAadAXRklehweUeayR3y92v1UWHj28lppfHSDGBj1kY+eX3SxwHIqAox55KZD46Qx5262+BK
dUNLTMrN50Y5CSpi9wXRukBFe7dIwxmEjYR2U9iezqan1ixsWpNYhD3IKLDZNRAUuF3aIkoNl8pS
4cx6vmZ+EZiU1bu2+VmCujAvpyq7Mf3WmPtzigh3c18Zr5j1xR+oJYAN9GA2UO2uSLOl9Pk+uL10
9YjqUWxeobYwmadO6unEc0R//FWoMgrQNLm6PnWarXUDKJnYU96Q+jN5Xd+cm/4gqVoO50Hc3MSa
1PeJ5gJtbx0Je7U8L/FFRVP8tZ+SOpccFkuoSG0EMXljjVtvxan+mNziVW2RtSImbrFfSSmnPvP4
+T2iHywpapRev0uRX6dWlkofMOE3jyTQ/Jw/Cd4TntdZRGhgiqRvkOOSoU4sN7OHaJqJYC4Kvxjj
IfVSWfpq3udIch7Bws/HhUjdyUOxk7sYhyr3yDhwrOi8h+2RzcYNzqMJ4wwnl5v3RLb88zrj4TYr
G1eXt53Yhd4SFSlkfBloMlxNydO0UBO0+72Pa+uaVudboJz8oWMWzRPxGrRYkR6ZQkscQJ/8fUPX
qp+Wv+5U1N8q2bUQmdTFd37WsOLw+YQ1K909A8hoxDErkEp/6ibKKvFk1GhedvW8WjuQ4wdJs7ex
8IkbddPOUAp07pRvAnN2NBb6S2//c/FKq5ipKYs3PqO0wFLH9wG1gR/8IOoLt7qBdg3k/L6+kM5X
HHi0Y6ObvhN7Hs3j61bdgDaxSyO+W+4/Wc7vOs+nnpZiXpZiij9MWcGuwmLhmUAYzpK6gSeLsXcc
TvvAn6brFHi4GcXgUFSyBov6cJFzbpzYTxxPjTxwwP1TyRECaFqR9K3GGobVUv+Mg5527WU3lCp+
Xr+N5LdEvGgmT2YJ3J5MR3MWkz6JjrFY4zughcZSFcDNIknNEYKsQdO0f9mT12UMitNaVvUb6qPo
6vkyQISOhIFAdG7LMuRmo1DC3L2rj2OGP9RVUY+a++E+2stmfdIi+u2SMIjcrJHQocRvIIQgwyUr
pRu0ioQ0RpnvpRs0cRdzKLuJc4Fp/SdkQqJr4Af6CO8DONhDYsqHO2GMKeF49wReewpgX9FeiSSl
RUQ7W3f8q/CEa7u0P9/pY/1wzNbjA/Mo9ABUdAZP2i/3urslmArZj2ADrwd0y4DJVNFrZr58BWsU
F9UbJE3lt3X2qUYgTXHR/eg9NEA4SqCnEdGHqISbFhsYbQDt2gMHjsH1RVHPsMQVx57vGaELG9/5
H1JaE8MnOUTwGtq9PEU9WJtVjaWmijdX9nUMB2K4nTDMmphSsprGQaFTC9KrULNWMKm8s6XTKRso
i3FBb7fwSd2KafgykjfJHwLQ4pn3kcx4eDl32aI4uZinIDcD42N75xBNrfma9igQ6x1LBDTIaqSe
6k7go5kWN2bEdjfBHAE5M9ibMHit6HwPrXFirXS+/kEQ8Wrfr6fY24duj504TWeHaL1Vk04wASXg
v17rTtCRK8FeYZxjXg1YRLSlUcSZQHxkhrQXIuNY5aICEtVAGwZpNw2sVM1j7lWlOG12upWaU9L+
Op/Wf4894xUm+DFB5gEYv2yIAJJAmtfW1/d3v8mjrHJmP7sDmkd5FRgS6wyOHi3MXVPZq/t3v76I
bYi/AMTQq+8Rj/07N+lCvxz8mDSqp5XhiXnDZQzlfgq4Ye5lzZ2cgeZt1jZclyGRhB+eCy2OKzN9
V68l133CB4cnpw+MP9L4pV2bI/2dnKomiojnZrhO+JdHlzuRplZK2+O6xbBH1I9I26iIOOLkBobi
bjCHB8mZie2+H8rVQNGzLIBgXcq7/kI7IO9iPfTR3Hhlib8rZnnFXZWDep3w4zQWjWJbneObiUiY
zWPqWrVjEUfouxBlvr0mvVMypr/dSei4yMlfS5bWyZ8vV9rAJUeA0a0A/JEgG9GlAxOgtGUcKcJ3
clolNyAFe2469ihgRxu/LmJ1m7lKpP+aJXVyDTJRqazok0XYiXUF0qXpZxQUoTG3CQUxBoFRM4TN
mcffhTny6Ry4WFxTZ9x3fU8F3MSaQXMU7VLolhRcH2f66nyR43ZXJNbPOpCrt4pY+yyfUhzz4Z4j
0FuIldfkBbkkxrmUTxU6t3d8/g2pwGiS7wU2LkApIxaClUrnXUgLnbYscnT8bZ2fRiid5apJJS8M
ob7jS/SyiIw4rEisejSa2iSxWS2IjZ00/cWbg0SNE286m+MWEgF3rNZyjRDK01fJHXOBdywJgqYF
vibKcDD18Jo41BOjiFRq77EywUm6u84Aifd7oyeMoKW2npHWIGuFmMV6u8ee4jriy3zol1H8BMJs
G7N6Hc1vNonNET4nBNqY/6JOzsXej5vrqsDGnPjt4TfaGhdyerZqa1W8NODbZBNq4f9ar0dQBvha
FsYLl2pQLFBLroTlro0/9zkrnCRrWfjUYZ2AQcpAibDzcefVwD9nHfSFJHoJav+5kuNMD8sWt1OP
jt94QTEybrC0KjYjyNoDpJUZON6Tgs7NZN+xbp7RfeAkTzZi2+c88eKyzPGGDR80dVm8AokVhSal
Hr1z9QjK7cw0vNpdA7xiFyaR0aTWx5m3ZdOtCR8Z+RGsC6zqaJQDNmJWw7HUR7ObnX0xCNLkUou+
llhQl/e45Sn/6I+AbTFBamJxgNWiuM6jGp1PTe1k6OTowbXeIXSW+vepmyypRXNXLOxplU0RoBhu
9EH7E+2OlPPa0QfhA+Qj+Qkoz7KavAnhBAatyQ01pYQ8O8hPvOnyM0HOkuhRyDOLGe/NNqC9YNXT
QcXAO0I8d6nROERF8wofNS2GSjuSpvjn8USQNmNu0mN7YJOcufbBIH53Y2k23Tw/FllvIDhh7V17
xOnKItPeGCC+DtP3woc4HoVZ6kL4rRkz+01sfH8pKSdQNqQPn2brrF2WBWjlowLYWnni0SrMJrnF
rrxpKhpngMoyeygvEh3vfxqwGPuNUArR7jm51eoJzQaHdk8F4j0fgt3Fmea6MeyLwptDy6IJoskm
TIJeM6uPX0Lw7CzsrmNyDdzu097YdmaxxKEscE+mdlC03ej85slV9nHlFDsz+1VZzvogJYS4oKTl
yGlL8JhhVAvHVNDI/okVqrB2PJOJJj/GkvMnxuHiEm9YM37OB+jy/ziJe2jidYv4ltsTWfL6yBY5
YgUch5wbx7CxXA0K/zH+G9NtXC6Sit6W+YUyrNq29emxmMwOi/BERyChT5pFlmpOiXJ1vQVL9Ba4
TQC0QlX3+oe2guNGjwEkHtFWlzJyzw8bWwJ5BvP2Zy9+rr9Fz6vydqpmawAGU2E/G6Vzx4wJhVNl
zni50unQj3OgDvwDyugyRcdGv5dj+zzKd4XsVl78wwUorHyJvaE9u6aWe44s9AaPu/a88jBxe0GA
imKPU7v7S0eW5XHeaFkIDfTiRxGkdIaa9RrtcVlycjIeogT4ldXDNeLaOoI0sr83lp5mRVKxINGp
/cGKVhHs9eAAcxpiZbpiWdkAE20gcvk55a9wGUfllaTChlc9JTodHksvROMTy5v7lZkLPbYfqyMo
PRYBB37eiFH7Nl2GGcKjWsHyzDM+EzGpPwzWQoHSdMRtdSJM/3crO8ph6hHNk5vnFnwdk2jr7sCe
/zXCyjSpZw/TE/PxA7ew1guobfSYbR1OajF89Fuiy8d72ZBKVBFpNiVmTfg0Fh0pW8G+ARLcqPAZ
Y39L9Ad7aN0oE4nNvF2uWt+1hKR6NIBmC6vnfVkdvJSjAq1jxK266XTIfO0eb/Ms/YAplX84/gjz
163qvdNJ0uryp0GCXPcPzqDBJo1+9fEM2Uox1RrOcjJcILBbOF/6Qeh6IWkiil7KmMsH1Eh/X3c0
3xZh4gZvT9F4VsIGmYirQl5eAM2tb9WK8FWfVp7NpAT9kTOpP/9qVZOO4m0RTB9nwvpY2hdhk8Wl
dg+QNgBc9RLYM19MTzXZsTfY2v7GyL3WT/Ulp1KHId8pFa2M96QMUTeqYts3IdLZpcDWuBJXHrEq
eBdSo95pwM9jQ2Fd5htySaTdCfbvAHpqQfXfOidscm0w41lN+/7kJbq0wDcmNKEfW4DbXtowNgMM
VCK9Cp6Yb+UjLGnK/jNp3XQkuF7GCqZDAX4Zch5NlvdecpCo5DeSmhVzEvLIYNI4rPxKpYxnUMGP
zGV448999CYJ3bwaXUJryN9bOuO80NI1I608UKpqEu7asoSPkm5ogZH5sYIgRX1dgCjkPpwcwFBv
/HXTE5opzbRc1erwROHWanGiERrCmEiMCe3dOqwtEgVA9tFOrWU4dosRQfBD28+tuWzp+VdbONtv
WOpLwm7ICzZNVWr85ULzAjMTLcgcpY5bRM6BcJ+4Q/1BiIw2BdLPwCFPsFpnnVFOtQm88KFxZi9m
EWypO70deC+r8hs2bzOuH37b27RMB3x4ENGdhRaHJkA78tCtGb4OZzANInZXIU2lBgrxCuVrmD/L
SD9UNfq/k+xUuKvYVke42Zu5qLmzkV3b8QBc+5y6Oav0QTZDMSJeRKKpv32eo0gCLCFrew8Y41DH
foy9a9i0pGX8qgYR8Wr8w2B9Cnk8MTpxoUp2PGWRr8Sd1HRUpsNJ2DnKPcaQY/J8mX8zIvNmyMMZ
xVb/o55QbRWQCBmrs66rGSiz/cJGGBk1WLEPYjrFY2AgvL7Cfn6cHLh4O/R6F0/Na3ISaIhwolqX
tkJ14nO5oupjWH7+dG+aqe8RPy+7FH6ih+/rx5rV6T3o57WnSzk7OTJGHyyeE7EbLvjUqjWv7bTg
YASW+L9zlayrLKGOTf54ioLs2HjMMJkrqiSXY/Bi60bgtgIxo9W9ZOunMCyqOYBj8zvcaYXYG3Jw
M5UMVgxU3xtmOgZ8cMKE4gDh20zJl3vhFEpnylBae2KS4kYLEc16pkyNP8NruoFlfIYNwMeV7+8s
tz3O7ERL8advCzD+KT3YKJ1IbZoRlS86rL8soXfyRMcXYxz5gbxTvn7hdoqMs+DE6e0DRhLpOilo
sCvC8schdHdArKJPpPuG/l+/CJuLbYGCaU0l90iaNp64wWRmbdXX27SlFHk8Hdp71Hji31JE315I
lTp9kbCUHi0X4dlbhQI9d1K/h5Vp1pPCenRnRgeLmzbkRlHMj5Yle1LHmRlJ7T119FWERpSSTFVG
D/xSND7UgclZsluwp9jnOr4mZ/Zg9DiLKhv2DjSlAo6m2r6BvoYBChfaFsgE8G0mq+VS93xOEeiy
4DCZhFzRHMpLcHK5TVGm/1gUgdCg34nqG6vDUyiR51BC+GmlqeJYcjgw7vwtflRO7tdRooxHpUS8
6gtlEjnKZm/rxK0IRiHzj25mYL/klUyzeG3AnXQCVOwm+BqxqM3FceP1DAkZCOCy/jL+ldu0xU6t
153UcjNYIHdUjsJKqRcHGOq2hwIyay7wOXmFgVWopJwPyTkqmXPGmRQf9ScBMs6TXtaG/jedLO1m
252KeCPlfKIdb5EAvC/MXvomMAadaM2HVjxv4PbPpYqb7y1CCWYq0jiW6Oo0ciFtR2n2uzaF5V+E
+md8HoifHlWLoPU0yxCJniSXsH3md0RNBM+2EwXnZVk5GsjQj9mrSEKuj6dmU5QaqAbOUDN+XQpF
f3IO6snFOAw9pZA2Z7+UqxqsG60f0URqjYKTYmSat03ULRDUG6mKcrA4wpWb1W+yimlces7IVGOG
dOH1jqQVBEUiYxvxf0hmi2KqPPdSyBYG6soEtgSRHxrp1JjqWmkgF+6unEls2vpBWtEeKCybpgKY
TBAaYlUfdNcN8CMB6+8T+M1kX5Xy3B8P2m5qNOMICv9D0j5sTXEgMMTgK/Js07+lj9bOaGymgJQZ
z2gMN5l/D47V0clTfp5xtQqii0BLLvL40be8/lvK7jLBCU1CuhX3EAek5E8kAd/w4G/rLQtD4bn2
JCHB2lCCSw1euSekdWy/V1gLCE3ONm+s4LSvXLXBUZTAhtgSAxxBQzwiaw4uruExSAlsgZoeom27
Z/TURymw6DERQsRDwabxaVn96U3GxR9ThIxRrShhIEKXvLmmepk1BcndwDFoo3bLamMXBQ1SJZf/
AXOPklWem/BjLIifFLb5xtAsqVZKQjkJhxWHhL4diyFwbrQBEEZB1WYdg1T5pdW+hOeGzzE1PpSo
1NHSsXK53CXirWMiDrKS+fdeQZ+i4H/6bUW27hAYgCrXXgaZRpGq/DWDwQzaDQsz3GDtGBhbT7op
T5bAfzrh+o02xsHY6zejmiQvetszIISY80gVe6bH6o1cruoCxXnl8k/fjZRS5s9wbo/+T/YHICGM
U8yHpQX1r4cERYWCip2Nl5BWpB9oW0rw4+C1xsiIFxgjMUdnRHb31GtL+1iX145SGZ3IQ2lAONDP
IXUSwymV1pXOBUOoloISx6VOe5/k9S8GXkMqPF9sIyxyn945oQviSamuMJtvWzYQcaVPKlRvpjh9
yjW7L8rXxCmRapGAoRclK6A/EdduS8aOmJuMGlt8lXJmp+X8Pqht74NCK6C2nQCawuFrfpHPGxk5
p5AxGLVtfvLos/LWHsyZAT5/hso4+lv4ibmD1Rc9Mwz+aBOq5AitqeLhJBklKgzyUtRIkQXbi4Bt
uxIRBoX6qCkBMrF4a7+uDJ40KcjddWIYISS2psOoWIsxayyhmVtjAPi35ZF5q24vhsmBZ6TP/DVi
U2mUU/7d/is4dm8EKbIYZdkgCnveHOlPDU7z01ZBFcz9hCwqF1Gs4F8Mj7u6vIjNgoyS1qDikJKZ
/AjS7yOAUicmfgAUYPFm9Nv4Z1TyJ3UjKKtSqAcvJKgDcmETu+IOOlLd46mVRLyGvwUNm3RVw8AX
FoJJh8iBLM49aiuH5HF2CJ7dyyPkggHdIZ22OmDrexTGF/xfi20zBANaZHheademE5UFdG1Z6Pdi
1uyFth6zYOO5bvpQl5aLr7ZkrrCAWnbGp0+7oBokHZopo3I6Ujc6VP/auIeEJ+SK1ZTGr3C6TnPh
SeIvtlxivMoJ7fS3ZuAngWXpA7k+Em5rjFaJS0ViyRrgtBe2GdYw4sUyc7Ki1pfvajyvFZiUAjCC
B1xXnZEXxVDvduveTcNe6VvqSbit82TTvvxR6DzEjxXOsyovSccGMADui3gEVc1vWKauuqkUAUyO
uH0GD0QWpEUN2ObmXH+s3sy325smVw4hNtaCn3e84yN8YnyEj3JYmvQE4qsXYsU0gKSv8Fnz0XWa
sGWmwXL1ELbK6BLIxFxPRsTEsbk37m3vnye53v2NdOGzFKQ8LVqN0bj8xKqxKyvX0Jo5sMUVUfbP
eCAKAatfCqFgHgC0oSmJKOT50LftfwV4mqecULfF9z38EovSsMB1QIzuDwj+bN4+MvXGgRSJu0q/
iKbBaygkHEc0QvghI8fgF6NNCZDrjLKE7gg/W5V5GTo2oT+zp19VLjcwHSKgw5vE+T3Hmq5zQvbP
5g8OtS0P5jY+nbOwu5nuh5AeCfcpHQkhOGhAm4bM9MMp38RVsXOgo5IYz+8PjS8iTVdLJT/KZGiq
9pCSu9D7XxbIkiOL6e4orBxCz79+Fitj8xmQzFV8CooWso99Blrqs/OW8+Q3PGDg7Sa19qMsOqWh
SipUE2OiTa6f/aJWBaAOf5Kw636k4GM8pTxFTgdeBAaJ6LmVmxyuCcyth9a0oBPCUFv9Wxu5M7Dg
Dtp2xb29Lqn1D1ipBVlLnkNvizGab7kDzrRP1eXEogXd0cIuy+X1CWGuQ46NJ+duDrH/0tNE50X0
eVyplZZF7pwkrdK6ijqkFpP7talM/6CW9OlMhDUwieW7CdIkYwiSKti4zyv8FPPPkR4eA/XTnWoo
hgyigv/471289/kOcnpMSnFl3W26A0eXK5xuJGXxnDfGRfTGKTcqEjyuXycf9Zh/vPALmUKwC6NA
nqzTUxRIWVVrfTaKUtQrXx2sAs3J+RBZvDu61BiO5bnBDbSW9atmWp6ZSofGQo0b2LzqJ5FCCb8p
tieLbTg3rAOcmgbgjHkpPKVsoh7fatax3URfRRRj2jRc7RKRA7c1Pc7vDP15eMoZw0fKHzgVEbNw
JalwB9jOkFfCcYWQ+lcpu1UQLP+y6dj1HrUd3gbJyVkv2y97m08f+qeeaQSvsMEhMmVpvpr5qTMA
ev49tDHx37aoBiXTNrZUVoIBJNkY+pWXosV27Hry5/HO2SidZTmbUuyUbUMrASaWvxmu7CMC/dhx
3rwyCnyDbUY7Uz/ZjPKDcfxUzwXEbJBq/Yfk0dGUgWwZv5c8Led/hrO6Vc2pGEXKxWCazorc3gS+
cPWE9jElJXAMYX13xFmCVJCxG/n5a9aHk0ZswEK1AOnv6EtFxlmG7CURwyDF+iFi+GvbtcIEg6CR
oye7o9N0YjNlUvo27B0oIfcSPXXCnef5cSp/QQxmm+UXJ1gVst4Ekc1tllwxPyI0zTSppMK8HR7E
w7VPYRQVPMZbV/wuc3dQ54p9ldg3TPwIkFqjZFJY1xwk5ICkIaHHNjfWHc6U/jt0uMbksMBcTHZk
JMZZDp05p1Nez+xRpDexUyj9rAOnut4cIsqzxz3t3PXtMvVhWZCQVZSBm4SvyK/ki+T+jYVYWAO8
HaSfr0rr3XgqjyrORpZK6byc4JNzXi617fwPPCjD8EPKj8AUIdNR76iUjbboPFsYovO0gt5yi6Gp
p+cVlIqOm62DEgYbIY+naadHHdPJ+EO8Xk/OTdcZyC1lp2s37mtBZLZ43PbshnLBpRgnp6XJp7yr
+5AK6uebGKBBHnVGpxe+rZuAijv1f4IjupqjoWdgPzLV4GppoW6evU0iQkKrjK5mrzZtijVokbAs
jaJvjHXDl8OVdiZNDbR+GzGr1R72mfanr3yqwIsfWS4dxdgGa7cNRYHwhfuzs+dPw0NKR3VFQZQN
eF3WXzjmuatDjQ3X4g7PtENGcGe+9Fip/q69LJ8wjADgYTY7q+PgzgIzOrFX+KX3lCxTnIYc8+HC
UzQS5Nan4IAKOW3CDwCEqsg/WIOeSfTqsChLOoPDSwN7pnJLJXAgIPjKVWLZQMMuwzKyfWNCs/NW
fSo7OneizbyTLtvBVFMLIG/RQDdu4M643mjQGePtjJ4FnX+8RyE63d0FaCaYAcN4slp19ctauTQA
wqiwXN0c0RPRSbny5zsEHwzqZ5/40Xk5BJVcgXmLWodWf8Q84M4kZrBL/6GLzcp9+WA183V4Kyno
vVTD+sezD+OnzzwzqsSxhAuGLJfNgoIx2+jgU3dyYTBCUpM/C2nXZkWV/q38NzSuiooVu8YIn3oE
CM5AuwPUriK4mBfoMpYrtLxK4USnT4LKefSVX9ef7imtxFwssYS5JqvjPS4mK2E37XKAKpXjAzVz
kbl0zxaXz58562Gqa+VMKW2QlgRliy2xFoVXQNqVvAS2XEqIOjksBoBykSjkA4wwvWfpDStJOJ9I
zUb7ask6/6Fo0w2PVP+P1uno2zgFxHFd+rmvDPrWD0hKv+SAqqSPptoYOT2/zd0a+ioc2DsyCMzG
wEdzxThRD8gcVfep7wClRCHgPX9lxv5Ov+SqpWd7zFTuStpFW4gH6aJUXiwEdo+sk6kjF8I7NPHX
GwFwFvO81CMfPRqADGCrhmdFhLLWv+gdop5c/igvEaTTT4k5pOIzv2FqKWibWDssSHXTW0VNQd+C
oV4HrjXw5NgScULI3qnjEeTaEs/EOo1Zsq0DId+iIOpUxY4rCdKtz2UXy7UxJHHq/ERxvjtwzCbn
wfyT7U14cBipvLTEl2tZ7ktmMPm4U/ZKXWnMFcz9EciF55Z5Kw9izFTQZm0Ms/BIoUOKjMHgcOOC
d1+K/Yy2KYylWE0CCmmBTH7LHyZp3T2QRN8N6tH49bKcwqcExPvIrUF2pOBtVCILpxXDHXyn8uRe
aFJpsDQJd1JE4ET5kvt2DvUlb44cAQmFuqA2tIINGj3GO4+31UNJAo6BIawvsFI8lk1eV4HaKbLC
IrnYBzR1Vo2ATF3fLBc6NHxDs+ns6pGjWksN3nRnPEqoxuztndnH0Tn4U1Eehm9ks+uSTbkj+8d7
uwFJO4nAl/eipQhsuXB1YmWI9HPy6uQQDAVMOSjFhLwvOMOvAMQHYxTIQQ1nEe4lUbsUMXg574Qg
ZDFHhoP936PG5k7LVb3BGWGLr8PZ5XdOh+992+ki2O6QaanW7lAq/xRm7jpeU0xo0PpEdcHp9SAO
Umyof505V8k0FYO5jHYigoRGzIRZqnUAL9mLjF4ohN3rWSlXLzIrcckN+RIG9mjXLJfoXwbjQxJ8
ZD86FEkNVyFXhxcvr003tiZmctGF+/gxCNMMbqaJFo1Mt2vH2CKS7NBPh3U8/jTCyuVjZweGp3C1
d3RpbP9eXag5gb/smnHUuHIVAHR/rCYzvmtoicloz/1pLYw6O7rmL95jbNLfWFSeAlQNoDp2rAc0
NtZ6NpbhIDbEOvbg+6JnyDAwGUSjqxOE17dITvkIMk/P9tBGUDyRGX/XYPTijwx9gX4r41OCOlKt
05TPWrW2Gd26Fs1w2/rD+GWBO4kmCwOmDthX/scIhFYthGIX9us/r7NtyeEcHDi4RqdngE25nE/Q
ZosRhlTLmU0PG9ej7UcRfyKim6XzI70MGYr2xo8NCAerpa7JfxkRGZf/eV46O/BXO7TBG4ciW4TE
EOMBQSea5E+YNxK+pxe3JbLmbmP+zMojEqG2/7pAz79I5JCi4SxVhymikqACQ9mZeBzAdP2ahdDM
/a6YHNyJiPTHJwwuQigp9tbGOlT9tLv431AOKRDCBqP6/1/mLqlTbtLfkYU/vxOl+yZlYVZ1dAbH
4szgydZ2QiwfoxpZnlpmvza08+pGAww3dtGkyBDV4tGyHU/o60iVWx9iRm3Y39UapvfVkGVZZrJ9
b+E2LWV3/zP+UpVE12tAtGJ96aeURuGWLCYDS4kd7qa6latUHn5zhbbsH5jijNgsacTCM2609HN+
pmDTxtbu7NRAr+qPcToCd+E3thFRFdXnfEhWlKaA4C6j4Fia76pAGUk4B0c9ZbJcluKUKS/O7UXt
4md+3WgfcP3/fjXjOUgyLiMgOSDK6saQ7bn0jbVAKaItIO39mFsLrIsjOhBULLeYwe1RhSNtT8W+
youdCvuMIRvTjG5pURsqRq2izXngPXVAjaoHRwVbLTNwaarcNs8ROWFfcrC5PQS3KfvvbsUppFx0
xt5iajCicdEHipMuw25JlJ5MpQPSv0CWWveMd+QjWKfxKZKfwp93Z49jWAd0tPxmxYT5GPRwGVyf
kHWlPUR3OWzQBhfpYS6iEIyNDLoM/AhF1EI1BfQhCUiY2uUIMEyjxVqoZWefEOR7R+WbKpgqM7SE
OHAJbll9oHhsW/rIzJf7JmoDN8eDbSWMcnU59aguw6JtZdyGE3ryCqT/pUB0gMPZ0K2ZcBNOQRYf
p1sMVkf36/qcQwjnTGdsZakYP5+yylSjU7kKk0fnb+WxFfMdYIUYl/VBOBYl4bL5OEVUb+xf6NWG
Q18dPEYsEfBe7WcGconFAZ1y5XKo/wF5ytHCGNY/U6hgGiEZQMCPF/WNx3/YmXoWwfklu7tsAHfH
xhmnU8ebzevXWOxZY1DfqSsspMAUgLJGfvowlWpE1u3cqvdhL+yUy00Dwqn0zspP2BIB8MdKLfp5
67E39+kT7jYXfCcUBvR8cv4loKXCgGjGWHmTx0Q5EQHCHzQAVUjBlYgh5NvtjlmFdvq/4h7w9Pm/
v9W/Ta2wIKb7RSIdGsA5WGQTzwXamY2v6eWtGf8ogSUfqYPu0uKgP+/agrvU+JBpJ/+hpvtzMYqu
mobeQfPJTXUMrkMnzYEJqBnv4rQ+gKXqRECsdpU5tiR2KqLgEWqJoT5bNrZr/ZMPdKnoVoiAbHB8
D99ahR/NLH2U04167xlZehYKf/+MDULsNMvCKZfvYmCOZ69k2Dqgsbyi8mgp3HqfEoKDeb2/jm66
LsEFayktij5UipyAvmPJsmy4F0cN6XGFriwtfDYPR3CW5oPTv+p5EWzDGRKCy8kioEuSBr6PXeEC
BZmzaH66bEyGqG57svCn3J4vMteBtmOAjSTlzlS/GO1LaPPdZvJlq6CdpdS58Xb/bQ6gsJa4yunf
sespyvwIWcz97SU8yfa0MXQxrCrKnQ6buM1NLSyOoA/cw+oIFAPO+4pxNvkyl1+Ips+ChAXSLiAe
A6xghlV2U2FzpB5EfHqTuzVJw7KYnd5NCZ70/OVuhm2gGQL6LUVFshwHi9vz14axFzdjiw4ceDA3
y74Mmqfc13iM9C5gUtNYDkZe8PXgXieL44EPNRxDgTC71QUSj++R1J3S4fnIHqUhk1W5dF4DvdNA
T41ZwWetdQ4dRC26V6mgHnCXHz9fMT/ThEJSzjGlf/5K94JFunPsaZROHEjFCIF1ejIL5iX3AQNm
DPJk6ZLkiPDUEAj5vNRGcDxMeOFuwCD5738SZ7LwnQ9GSJ6TQwnl1nRW3U3zt5GXd0cFhUlEw9AX
XUoCca8cFxm5AN8h9ZHBz3Sflhq9p2u0WQqJgvYLWCo9oferF6xflS1DdH6LPJk0S42d9oawffUx
MyKYLzzNbG1ArSqqyJiTRISRRhue76/0tOOc+PC3moh3TGf8d9MX9bidijBXGwamTz6KtD2kw5Ib
XujROwAAU+qOhqGikDUFLbUuJB3yQeXM2ENOvExQ3JTbdJm8T5afow+f3TJTnI82sUQ6ktRu/6M7
CuldgrwsNbyYqwkQnnhNZ5FFj/rXdPATgJiwt0MHRp5mEmTbPEc6iqbB3rIkcAqclL4ZZEPjzDC8
R5k1Aa2onW0u0DhzT+7hvlPSNkEQDjIKooLs0RsgDeq4QlQ1DlCx1cGRsWH6ZIMyw2d5X702FiDv
Xy9MNPfqTbbpIi1KT1JW11BJ6vSDTT20ppbZt+bkCDY3ill6p7wJXgo6uKfqmbn7ZnMuamI16s7O
LJFSi7sjrufhvezQttlRIwQBWgJ6LhvDuzOB6UaQhSW8AlKiuUUCGV83CudXAOxE6AMRKukj9GwD
rSIOkrOluYvf48lxhqFY17IgrNDu6Tfgyrb4H64TF+C0oARgPNRKSKF2pZAzBlPDxzECLFjSo+1s
qjbyMvYRyF2jR4NaEMCpFU4x+FFCMbTV3wl9oWYzyU7wJ4NQBVJKGAl0LebBUOK2AuDh/q1Xlc0D
2kwo1W5NzTYq0nTHWyDfk84BefIX2hnBdjYh0xWhqZ2bp9JG743prlg9uGTpCzpo/wXp8J7U2ZMS
GeWY7YVtXXoXi/RoG6rEailk99RQIljfdD70aR/atxR0DPua2CiRqysO2BGRmZePGB2yzch2Z8I4
dNnzlrqL5ke23N0IdCcEQR9eDam1OGH7AkB8TeGiy4RBlRIadTtP1f+R4R5oHVrJg/4DYq6AwmnV
nh8lGWe3A//Cy4oxxAbumFVLBlVntz3bItuKzKUyLM3iziSC04DoWYiLPiuEGhcD5EA3yrLyIrBL
vmlsG/ZHvPA03iSiP9uSQ0wUsnVBD6M+QneCsMiK+TRhkwhMi9dPH2653QuQ1nGiO/E7RVXBEHmV
vDD7iJsLL2SmpmJGsRbTIgXzZni/5RXGcetlTJyq+tcNfc55Z/vGIWqKN4ilAOieTMPKH+Mk/jC4
nEk/fiLPWccm2XTkulV3HwSz6IVmEWNXdZEeqaGK+EdMAzEz4KJSHHoZRxwJ4B3Xve1i4RgFGCn+
nwiY4p6zscskNgSqsPsLg8FYTesVdKYIzKbZWhAvwz8fWgPMMu/L2hH2UGVJ6B+t/auNpxOhogZz
PQmWFGyvUE3w75v3UcMKc4zF0+1lLZZxTVijQ+Bm7fnQzIaqeHEMYeFFevsy92zuw0HLWwhmrV1+
83KreobHJtmH6aLfCAgNvAHDF89t+pFLP4UMBbxi+5kSo/QLrKEmyFccUV88mTDKO2Bz3Mp1NfMz
EH6wrJ6u4AO1GaFsBtD0j2TGc1g/0KML7x+z/D7pTOnZTu4cYdzNUg4ur5MDqEvu/PCncVQJBYqL
44gsg3GbvDocN8Y/gcxdYm9jniEzc75bFl8YGFPaZLpGCKGLXd1ioz+YMl8+/88xHDrnpgUsQNCc
CyUVQNTYdrY6lB7JJqy+QtzVKs80u/dXVa4wYFl6FgKjg+4P0lCHvkPa3UMdbNkJjt4JrqAk8yJX
sO77Gbez8bacTfH/u91A8hG7niqcW4KMm0mZimsiRgyw2gc4Oiq2dKtoZ1ELdVRWXY5aS74ICdxj
J+/KOb+8B5M8rPLUNKUXpPh6DYaNJ3WU032CcEYv/hVjMXo9OjtKgeyNTbPFvoke5CYMVJSUidMU
AtOudp/HAs0L0D1rMkqaqK9MWm6M+nI1oMqqobmQvycT5uVUm490c1YVfMRHAgjJNGZreokiddB0
tv8DFm91+/hvWMBQcNPasgRno0uEciWAQ9fdqdPHsome/AypRwrIJcKyltBv8uauxbLjPNiKqRVS
/x+qhK49HIy7q2zR4ArAEuSa9BDh3wcf77DkL4ZqzKoHf9CHbkrwhpERCuC6Tef1dLDX4KJzAQ0c
AKfOnEsvu3swsd9uR5HWqvwASZjnJN9mONNNjDBc2SW+vDM6KAXY+h0pHMYBi8TTSeoxRZ7rEaEz
vu2MQDDNOT/wsqJ4VEyoj06xB//r7PLZd6osBMAx2TRHKT4ABdISzzdLZMjsJhbb4x0mNlGSUpWX
mGBmKhLU4T9fZHiZ6zLZnMIlxMWLtU+RalDl43ZHqS7dO/MIFWAcmNL5owZ/Wp32y2U8nv7fe7xG
6DoxrYUgRiy1NURNJPOfRAC9ZEEMpooOqZSlNhW6HyWxmPqewDeaYLXTiGo+cqeI5Ho5hzrqxHBf
Es9cNwpV5jac+JdAtUELds9zDp52QNJ1DeOcq7seIi0KcCIB/5St0+Uebwomf5Fveajl+yP7jAxa
KIjlYJL7iUf576H1JhDdF/3xZg/BMdSeN+MJwD7BPW3RGTS0nKdC8LZGSfqNcKedPavB1WKCUOAe
LejMluHzwUPW89WyvSFMYMeJViqJ4SQ46SOmcyCryGoRiylU3oHkpb6kRaHoBFLEYdsaJ/6qwUdn
Ye4pNl5KTPRLP9Aw5OLbxIyOY97hPHWn+OulDMpq6qNvJObWRN2q7Sw0rUZryUTqP7naCWh8jKAW
zrIxzZbu4Vg09KbGBFgk0OrmzaREXLSh7L35zI8kcZm51AwsN21plivU3JUXtAygBq+aTQ0/s81I
o8tp0YA5hxWIm1gaUlJ77mT9YQ/muqVkt0J61Webpi7VIJ0giGFnZBOjNkPc66tM1O9wfDtziiCw
+mKc8EmsO48Dp3QdifwF8QXIZLYtZu5rFFDij2JDNWYWeBMFN7Ig7cUVXntclQPclPLcd1U2naZg
gZWhFGU+Vhk6+seE6Z3H62IyZXLGQoTNGsD57na7HQ5r/lB/jZl2xiHmkJRAVv5A7KtSLAC3ZAwg
I82ifTe4Vt/RdTU0jyx35A00JvkhLSR9SL9OpAxoDQrKGyH/5mumyM5Fim/aXUVze0Baskelxbtd
2jk0ra0loov66Pk1bXT9/g3HGMYlpfCvyG1iOLrQoB551qagAoMQZYKU9vx2wa8lePrsvaTTwu9V
bIHlkQ+86wGiYYyeHvWfFfiATfrdaT2XftYyytvgcMB/cwvYfEP0M0UG5QZ06DI4hFpm6xLbxuxF
uIWBSyP8Oa4dCdaHirik3uye/IzmbJCIjZcTazHW5sLxZXjxQ6O1Atmz0HYzQH6B9ixdsG+qh2g+
xYtKddoQXnMSAiA++ZVUfZSIzqk7pfk4ELLysmT8S/JjoTKwQUuTzM2XF1rqVHkbxvemnb+B9Ps5
fHRMSw7Ghif0wbv3zwb1HyX8MFt0Q+HPiRmntYh3ybCNj3BN+cUFZHrD7iQ6ILcTgvL3HTB/Age5
zheRe1GMMPj9yiqwpcXJ7aoyVs/mYRE04+vAjpoWKxgGBYjfOoSpKuu1d7Gg3WZX7WoTQerbJ3+2
+YVkzABGgXl2bvWLYtt79HMeCFD0JLXJsaHQ/drGGiHxyNAH3MaWFEgf6Y+PuXLMpRt8d9g/8PMj
iGdx81rWTh0wIj5co/el+Ymis7Bp+Fo+BQZxU7pnKNPAbFrqhSTWnzVLiWEHGr/oOjp09Bfukq7u
WEgPVJqZy0Cu27giK2j18nyWYwml39JiSr31uM9dQ/dYvLeidx3lXsDoEQsAIFpjTPsr9nO1Mwtw
V2RZpFp11897ukoZxeZqNJjlYBEB3Rqn92HmXT2BJzQJU7C4edSvF34mQUkQUdWdOAW5d1Kgin2W
k2NeElGRn2WiAuhIhjfKI3iVIHzw9x3TEWXd3Yzg09Fh0aCEDgMS2kSgBSm2Ccihf8/gs5qYWFGA
2geNXDs6RaNds99JZnVH1HvQLwrxTjzb84GjwiVINI9LjnVyn+Cl5IpYaW0DopzL9upJUr/FIj1R
QHesGMTQ3eEowwHrPcA4bC3V4h6hatxsvvAKCnJCzGB6n4bKntcYo5y2uaAz/3DT3TsBtFahpP+Y
qO5gZ2tqXCdrs/6y/QUPTnhNXedVgdw3XbXcJzLJDmq7D9TIVeYxqtSBLTRh+61jIZWeHSaitNJx
8OtPhP33JRwHiIaQnvU02TXecM/VuaSAoeAxgOLODt+fLYEneEUxm/sFufXQID5bL7k4CcMIifPB
Aer/UVVVhebR7VoZ+Exr9Mzkjf0Dr/VWYbyVr5YrvkUbzwn1HTcMRGRNOQ67EwS0UjQQ7vtYyZSN
P4Di+j49KwBdlVBL14CAatzLinSlGXyYksDvezpIJsxGLfOhkxcdAhermthTh7+gad+7v1A9pj1/
oPDy+FZapeIDaXtOYDiWDhD3ChlB88NekjyQmKezC73dAK8qsO6FHpagzmZLJRIQ83Kh1OHBRqx9
CkfhBQQ+cPh7sl09mCvPnCGfQEU/DdpT2C/pi+aH74NEgbPjer0EEMTDH8uFOr+bKr2nmhn2Tc56
bLGX7dvxPJQ60MA89EfscOEA0FJNhJDb8+Ju+kya62Fm0jr9SEcFcbGt0nVwsNClH2YxiAmOTHZe
Vj13tZOP5XE154h4OafaXbydVW+HrQU/KeUI2fkNZPFr6UXDRpXtlIIUiyuUpSDeV6lKJX6q3Xgt
UuOhhG9Nv1tXQKbpF0V/bCrf72RqnV4fyopw2bjMrpO3rI4+4UUFDyELMAAx4rVE68fI93Y8p3OC
hWLOIioRXT2pI9a4/PQ6PITmhxyv8Ss9a1pdh5cyL1V1m86DLGk6BFAA6upYV4xqWtGIoGctNT0y
8HXWPQybsJXs16f/RcHLnwQWDg87ooZYeNrkmw0SHOBEegrc0uXEAvNS9ZntONCIsDJCWXb5LQue
km+bURJOl1EzCH/uQGjjajm1qKk3dIKuSP4Vh6W84YDZCNZsyqHzYcgwYLV/MY3DgSa8xcD9aci5
+LjEla9Cqp2ow73wRvlEIpbZ53kFhr88UyqIHEl9ay+H+GgWbDVdAEhA1C+47RnlFcODCWxsPqjq
CIePEZyby6Cte9oyn/uEybJnq2d1oJav+O2uOL7cOGJXIvLYoSmzQnpNZuGlCCWGDRxnKpHhNhcK
iohsQG50PkV6CTaP+u1V08RMvfcLFMJWFHuffWBT6eFUi26R1rlO0GyTHte3zux+udBZl4723UOG
xsMtbC7hgBwykbFKkD30ujaysjEyIruOuZeXYXDx9DRSHBEUrPwSIBGYk5t1MFfR7MwxCyaQAVcm
tbKPG30J86vi8yAtIyiShT3OmN7lnwcZovVaj1x3/3LAYdATRtfwWFj7VFxlEfk0qxP2KpDAdPWl
yVDvaGKin9mHuP9XnNlycYYYKWYwwPCOzsa+vIpnAyzSS4f2rsmxZAa7k9STDAUf16+RlK1wYbxr
oc1JKrUSqNsHKXX7NJ6V2EqlrZ6n6AfsO/9jpPA8gm/QiXp0LzmjBKoLGOl1fPvmXaIE4154O3Xq
XEAl4TvETe0fO1v5iIUqNP01cLaDRtd/6P9HihqjbTHqsnbjcvjHI+f6aWPUlnZWncwVwbU/+TpZ
8y9P+tZT/D/5OVMlVRKTcw/KC6H/iMNJER5HK4LRMmDPv/0+JVBeEMioS6u2jHTBmyv/pxUHkmLU
PP+zbG2Ftmuq2sftDTwAOkgH1XbbNk9+MfQCAYDKunGImsGroywkk7zu4pb9J0ZOplwYAVl8qZcs
njRWJR22uoN4GN/C2aUuyUZMAMvb1QmBwXhlVEriGeG7773N02/Ax/lrhAbQYKJFqV2QR5KADzNd
d6UNb1dGZsR1K0fmZJWSfNsmPesNQKzo9vPOQn4QqweXhamaVXb27ETTGXiloKjbGeMqnbfmKrgO
svX3IG3ZuxQ9elYWyx1wpZxbJ/1J0DpXqjobOwaIyagA293AbVt5SMMtWAfjZnd6FFJ3W1V7zzEk
vnSBC2i6c1FotnnrhVFbOZsh+ly01+Y34m+JNzFNZ2Biti/VXX7mmclvBxSd0FQAwA0pnZLnNzEu
jojy1G3J6MbcgqtvQYvOdKeyAH6yNHJmQpdTAEnU5BDCtQxpkEYYxG20sYY/VIWc3OUczLopyFuQ
k1IrrgcL1zXrvRyBXJCf8o0fcAJ4p0XblfCRyOedKwhfq9J9KTTQ+kot6+TaWubT3rhDjbr5uZNq
jtVPaKR2HtiQhIUlQyrHMGSMjASZYoh/351V50gWqfQWFRUEd1H0byVz3hyxk0JH5xq81C78FAqX
zAm3qh2Oz3kwSYO94dzl1rZpaCFEDkaiIG+LNe1rijUp6YXa+TqTVCsemC7LawtbPQ9OwZBqNRUq
vXft5Ty4Pu451F7qMrJMcLJKkHk0qHSNdRXu/l56aEO10Eb1KF1CLOrfxwB2UYGUpWx/zJ+e7AZg
IIz+8uOJld5CcKvnRVD3+j3+qnUhG+R3x+RlYcCSkYIR5Jxs+UYuXShUv+BhivUFhP4VmbuRAHUp
9Edbp9YSKcnNd8ndc92yzQUjQH69bNvkjAfbohoBoSP6s30dQN900V/yhjHlJ2bKm+tQu20LTYEE
C+hhvS2+BUkR4OJ0+DBegshGdTgxaAsdwoL69XlVabuVm8rv90f28tbcQ6KINNRIUMgXnlvzFTGx
zE0Tylx+tmRjzbbuRCpHswaYtp1c1BXBm4UpRZjBTEoTr3oulJTUrkDKZTR6czABYwkxkFhKTznR
bt5SGWysmp7VBaA2chWkcCxM8SYyKZ0KcTKFB6NkREmaiTu4UBZQKtkBlrMuWpyXjV5/U58iWVl0
vsgGGiTzYv9H8EfSRV2j2fttv/560JlW9gAN4hrX7pKyzSbBX9KL0GA5KNpxPF0UsFGh3eqNlRaT
55T8nDC/YQkneYs3vWWODR7kLP755VWPQSIyWb7AgCsC3OdioKk/7SRK8PPWZeaxSuXn4W3Dr9/8
F19HKJYNTgiC/rfV0TrDROwOL3lwg8S987dfYOfz3/RLM2TeFe2LvTeaRRame0C5kCzJOcUcHVTR
1Pb0PtODS5/X5dnnCOHtgukREZG7buJRYyZ4BlwUh04pXXm4xmyAuZ1+Q5PlnEMKGpjCrv+2VUif
0hp3uibixfyz7DiinfUj2bZOmfjS700Bh51A+7JbmK3TH4ztwGr2uyITS5WQzkvMCCHnoGXvQgon
mHBcc0qGMWKExcabeooa9U4XTugW20KP3DMPi9Gj0npa8QvasTDWjzYHI/QOtyzVO5XD15KZ/Q3l
i5JZ5FMZU+6cgVSnxJSm+nBvo+pFcNlLX2eY2/pKYnmyLjQ5XQVrx1A7fQbqB7azdP2UQrK1NfCs
ogffXjza1CeKFI6WM0HuO+mv60SwC9Wlw68n5FrYzvt2ZKtKRTaoaZDFFzHaizCwwEWJzE8KfdC7
UtAO6KUDAN4dod5ythf/CtE3YlypQBxMCUMAYI6xK4utiTwSTJg67XgbNOZWEmt89Jy3SbE0vAPp
O5CGnkLr4gCfAmjNS0itCbXuuRKZhJ2oHG5axrRk/pvrfi7kPiPHXklURFyLM0KEtY2B/3xFCs+T
2HVYBGv7PaxggjqAXT/Csg8ixNWu5prWPRUdQu6Tudy8K5YdS2ISC0G58y9P4YoiDuLRa7VAkAoG
lIzQq1mIot3RNrgvpd09Z4i6TJxfgaJqwvgDE7oyQgd7af9v2SVMrOYZcy8CiPor0lOnFny6RncP
Ld7EH73Rszl2hNAsfueuB9mII3sahnzCKls1wBata+GHvBZ5pFWTrByGyE4iRu3EAk048fb0Hpbx
sFCS6NbzbSEVNPNv+78fypk1LBCh24wZNHoywy2jE5E+E4KGPw+p77fUiex2wAAS9TfvCj/iZ0gN
Irc2dj8JlX3XrX8a/IybLWmjZj3HrHBP19fNsFoqK+pwH0JxwX2MAz7Fmoqjz+J7qPUDIq23XPkE
if9TmCFsHpx2L2aL0LXUA6WlZT1p/VsLY6wuoO3r7xzgMyDoUuZLn+PpAURTPlmVqvM3x7NhVBm/
o6qf4Ck5xtpVAkn7pRV7afTjsaEPXWUJb12b5XKkrRR3SyPEla8/9700tNrNSKQgFV8jOid97je4
ntasSObg0RpaJAlHx+4/kzFliyPkHVFshKHendc8B/wbdAzoNJWpNF7vrHoFYspAkUTGbDON6A0o
jGxV9RTCCTMj0WL/rcoQIB+TLRwrEuxORaXa4Zw7bvNdV8+Fxq4e/dxxKV94RFJeYiAxurJtN6QH
WiC1QFZvzcmZIJ2iQ8AjVpX0gw1TCFXRbvpEJgadXSLCo76u48X/53P7PYMgEbLf+BMGkek+dJHq
yl1HoPj+HF4WS7RN3Y6hgJE3yBoxwIOlQ978bwvc3bNbc/eH+1hEKxW6rgUdYSKdsmMf02HY61vY
QvX/wlQaDrah6mfNKW1j1dvSPkLxDMSLI7uwni+/V2puH416weaK/TUL9uR4vlrp6+8uqHF3GCJS
dMciS50wwmEH+bZe1OLsG+zIWYJ0XyzSbid4Ti7JQ6Z2YwfCjwQngbnpmtQmmbS2DocYebCJWkIe
Wcn037ZvRsHvSSuE0tLNnfSbodWhJ2lNjy2rByRPastcI+lesMsnaW8b2uv0FTAbUEQhm8dFtqgC
80npBanLWCVw42DrQ63DZfmJTOKNoG02gyUTPDGbsrnDa7JzkjwKA9UtmS7ZLEVCu0oDmbpvjHeJ
cHTYJnPcmwjN/o64uoKZxyY+NHZFK8eiyInkifd9w9eNlVb845fbkWdg3L85eN8ByddYcj3sUnzE
dohw+OUi/DtQcZ8itviSsMzoqWlpmOQv2lLMZMflyYcsmzx+0FsY6tP352i3dG41hPFyhX4eP/Yd
gk+tvxIY/iOJ9eXibB383CZuraGyRRu6yekN1Opjde+JRVkkmYwpRH3v9zdYrH3GucI7Zs7BC5Pb
X5R8oe1AKpN+LhXwtdptmoeqslZcfI/l3ZAb6n6oA5ATyPxoVeHwVG5eR7ymVw5TEG8z+YeAkeFS
frOXrlJyXaWR0MuHEdCbOmCa9xiaAJETrrYY61CKS/PzsZjfW8QAACamcOlxwAxWIIBZb1yThuR2
qGzf4grrP/b+zhP+rQoyP0Ztrt2tPYxK/KgyRKCeJPK/Xq3wUkv9C8itLIo7GnOGp43FKoaicPb7
iMcoFNLgsfg/bPn465ZBnAvytRyyXvfeEb5+huW2st0J7KqmxIWABxmbR4vZNziJGQOJz/IuTO7G
kmA2xkChzZvr4hsAkR9d1hHDj2y7gUoG5TWkPL1+rz8MSOOA8RDvVqDQfz4dsHXIq/ZaBFNkNoD6
B96zXcRV5M/DdYVN/O4LYbeynR7t4XioAmvhzJdKbw+dc2qVMvFX6kl3KM9qySuJxS3f0XVz/8et
6KJuE/rYfytZYu9MaJERTjbQz32T5zGFL6bWEUuktHJBVzApcAzSIhn6KzcF7UnHnrmpXtOgDQAz
vxdkQR8oeZJC34AanbgeF8J0w2A0DUlObKYu4HS3Y69C7UT/S0BC8wyAbl1FPuE7TbTRBa8c6n/5
YEn8UqZPSZsBhigskNlaOrDQ+TFnErF3arwjY2wySh12k7IAYnIMT9JvSteTACy3hguQOnwiZfIk
0O2Fih+QMPTKyqTJvZR9E4/XtTDRCMYeuPrSnnhitTwAOFluJZLQJ67i4iPYfuxrrrU3ki6MH31F
6Mztw5FcYtZzWAwG6jnouDUoNfsRdS1E5ljHf4eUuh2A47CQJLja9pq00bPO7bshHfypxAl+tqQQ
f3qyOG4jl10wBVWGVKvy/uL3RCDdEzRbWm9EtbRQ/+qHG9Lk/suf6M6UP+XyNm/aNvI5tq2IzQLl
WfrO+MBPrLWzaB9vK36QooKRaGKYxmSVQ36chdWYmDfbWx4ghcKFblJxo8QTGzBL1/ggrdCgLMjy
ZiH7fYYH9jF0z+9sSCuV8uu+fg9sIaKLyYI0EjfeW1sRDiXTwHOgMry1S/OQjA4zWU7SNr7zq3BI
Z3FI0i+dAUbDdolE+S+s0S3TaMu0eVSFvm4ofVAZPwkQXlcGVDHqa78+Lj425/VdrK1cmLb4oU3H
YrJ0qTHKdE9ESOZDU0SBzxzjsgSej7Yt6ToiNKwHSmkUyFVOkT0E/7xw1nG21jhLivmFwC5tz7jR
cvR8gSa34ZGBXjxuVplAj6E466cG/OUAn/QfcuJgYQkXezY7Irod73DD3Bwq7kBkaqVV7s5eTy50
zcMeqCSkj21uIHUYcuGRgjYXSoBNDDB3Ot6ZMy0Z1yF/UzMiA/azmEdZjDTMnir9C1NWnPyIJbqw
0U+FvunCT0EdZpZpQ3fkgWURMRQ+M1EgtPekbT9noVGEgKzs61FmEmHnThSE+JEbxEHsxehvqZjT
RDIggsMw1eUxTZdEOEfrvlzGgd0YW5pT0YNjcRpP0/ycAly6GQRqDNNlhm6mqWaKbZy48UXt3ejm
gLwuCez4eDR0TIRpw44oY/6rDdTudUNp7zVra2ClCf3bfYFuEJnQIZULUCOb/kI0xyQgsrl17rj3
ahPNrEJHvOAIGxobPxIBfA8Wz+SxyZR0t8Nce3yV3+nEJ+odDqA0xThBK4083ujiHQ8ZF3iIxTHe
wAQ9sv7wqVKwCyFLVw63kCgdEZGGkVCE0q4wdVn3Sz/o8MMRf8MKr9JtxxnUTcJcnqZ4ZKAoTZz3
oVNZBjBhA8OTS7T1CexOMLJHn4hfABYs/c6z/3EhdkOWsMzrtEclPKsXCGohFXQXKBHCy7npVinP
C0DWEYG5q3ko+94262FaHEXJqB+zonl+hAjxdb4P5Pjewx6RvR9XYsYmNKGPnB2+m7716GuX2TKz
vuROJ2DTVGOf0l3IKFLTmGjMijbZVHezyNFFv+wkya9/3bUp324uAbjnhPt1Zpn0YHaroBApBnSg
vrqulvCAnhESY3dBDoA5dB45lQf91woPJxiQCkQgWpbmpbZKbDhLiQtGQJ2tuk7/9EAJjP6eUPPx
stInbZzrVhTpviOltGtT09HdxlcwdwudcRPbfj/vheKA5yDNU1rRAWufK3TD0taC2M8c5gIeOVyN
jB0+pAWbl72bhExBY1giCCyNO9oAZdoRvSWCcqRjckuXLdrhM0Jrljr/Yw2nxaRCP+2VDoM3q64A
xls/60k3MT1yIdq2c+K00Iv4izplcaT/r9vPDC9Wm0RZUiQkWBXXMIJVLDbWdOh9dAj3teU/Qwqf
sPhn3L6yNif1090t+hwbqf/0+iqIdlKtQwhsa95UrOEO34jUlTIKa31X1em54pB8EWy7GBSAE7Ha
eO6MWfoMTxrQ8SOOtbom2pJE4TqNdIqpcUTQ95tmHfEadD7qGuDSuiaGPEd/6PFIaSzanEy3fC6I
iWPK7hbX6XCku5kFXpNJuJ7erhHFD48Yxq7tFKpMMXQfbwfOcL11q1MWZAmNZXJ79PPG1F6Dh+rv
qGxe8m/BDmkcmBsNGrntjaV8xwq2wUt8N1chVSdLIEyRplOKWw49y7rsY2jX4QZcYCQBkOuqKcBn
AH8BIAZIU0JhVh7+7hoJ7DPeRk5Ha/92buFiPClSyrauNJlyDIN8hKIOCb7klPIia+GNliOFjlqm
zsOIRAhCihA5Fs5TLylGdcPwj3kJd8Brhn8SG45GTS+NoNUSk9r5EbONLHx3XYKEcmmqDPsShnlu
ExH9xJBStNZA0SkCvpnYaTwRhT+vZThAb2/97at9ppw0B4rcMHGegSeOq9y8Oksukgqibe0+8WkE
rUJ7Mb12qssFgwS1xG4khoyHkGmuDTFq0n8NqZxYZeQJ9HFoQc3Z8Tlq4TcB8xOOWDTnlogwOKlp
UHpLpdTcQ98RAT0o84+DoCDZLotH0W+dcTD6pEUZ8OAwfaadlCcKHMV5Sv3eeQORLu76EyRtBuWj
bObG50zJ7JRka/7A6qvjrfNYj7Z6+qX2RqXbU20hRnCiWYJSTt04vefUpGOMhAqOYixgvMAbSvBL
fFhiOlvK4Tdz5ibnfsiu1nuN04OF7HmpB/K+mU34ljgC15DK5M+Jk2JQuZWDEYWnoqqaSN+buT5h
JfSPKxdHKjOdgU3S9VzmO/gG99J7uoMLVqrIB2hLpA4Qhwtti1qWX5pFosiZ4ed23kNGstDIOssy
1HmrzOp15n8u/YKuHlRKTkALv5Hh8lkezxYrSyxEfm2qGxgV3JmrBWgKk63o57ta8LIUECBIww8s
fEvluZPK7Ss7s/ZwhFveV8vnhCsdZjjnJ8/g+axz/eESS+WlQPW4fsg21gneCmZnZet4moNrmOA7
a9+2Z2+2zY64qr4+dPpu4hT0b/XmwimlnwleAOEoHCA7pQG6435N+uGy87eNZN6+2pDyv3lkroZg
AU+U7eutabYtq42iwAYxR8CnoOw53t6n53pTdAUNopTDMydDOW048tnkv/yCJa4+yJSYDVMWXU+J
o+vN57nlw2w3BnL2XhRTKn5L8Eh6pDs6hjhIgB74oWTeIrG6jAzgym7mvhtxnCgrUmXEoMYVe9ui
6HLmjxhsz1w9I15nEhlvOwRkSNWbWWbHJkkLlaqRSNH80LjXyEbjmQdUvFF/RfoaEo1Pe6k8759r
/6J1XmrNIaaFnRmGODjyjBl62NZV0I85dmuAA0xkKoh8rTvHnwZlGTM4NDB2iJocOZQ/NMounLFk
N95C9fdBT2R0Ay3N/tXYlW/FvVgP8JvgdB2GHp9sLmLbzTjqlLySzQ95CLcDooFnySFPVHyqLEm1
kMdxGAqBTsBC//OD+GPuMjr3eOUijRjRMRnt/Gceor8k6nz4vmRZPMQxKuJW6jSiIDy0XU7bwwHN
+MZK+gKgftbWX1E9iQ0D9Bh/J/A1N/rVulu1L7BiRtfUSDpeUxjJndAn7Pa/44ACazFvq+H8Qsvm
1+MbUPr2mGi7EAcSQNCWgYj5CkV1LPnZLbvwrU+6KUTkJhJn1y1E3rzfwW1wA4yCvJCc/LjpRuDy
TcG9c2z4MykHZA3ZuYLDHKTQlFncjQW9uZTr0CzCJenjqJGleQzscYCqdd0WV1lzKSjuTEOsPRSd
Yj5w3JJeSxP5Ng8Q82wisiUQ6pWWPCWYiNyM4NzHRxtf5CCLeqA+eMpmXLL6s3u2+kN+I5ghjYEb
hCIWSzLUI99S1rG/CK+k7D0IzRBrQffouioHbJTylt6y1Kfj1irp2UwP61Hot28mt03zWVTQzDlp
ctVaLqUAy8PF1scIuBhPmGvHNJRQJvdyFMH3+OO+C8zRwy2+y5ofkScd38DNK9xyXfc4gsZWfTOb
o5tTBwShfn8DTuPrC2/UIQC2foPPs9XTLKaIfZViyEDSOgGr15nREbxiFW8ICNXn+aETINs8l7yR
87VNx6DfzrVZC0wG7UHZptDzJHON6abYq4n/5yQY6blOsO0AjDJuL3ep8/PMfv4gOzqivunUQts7
rIZRHBWdyUd1Hn3hAOJI3JmpUPcG52l9J5qilvQ7RdHsBAlH/2mcLBQJ1SCAE6LpKshrP+Z2K6/r
D78rRXsVexUq9t/T0pLMN0wYd+3m6QSS+KoMk8WyfuHGIb++IZO0hEsYNSl5URBwJ72flyrCXV2+
hK3M+tQPh78HbFrZhvw+e7tcNl9SyJNGX/UVDnIp+gYCYgxEFhc8nJKatY1gXBp5+JA7+AOlCidY
rQvtuBb+Po/Df1mQ//kPjsqHVh9BImRAMvZoUGQsfVaXFCMGgAH5sKK7HjOChDRximRzIA/AxOrE
izn9JBWD4ZXi7TUXXfQcWMOrvC6pvaIpClWtSmFj1PRmUXqt2CbwQuNi6Sl7Hzo9LRq4zgYxIx7f
N9r1M1q6mEIfMlB318l2ggxcm6avSH+pHBYSIHywUyYnHvtJcj6cCJC9v1LFnM/ngfWFVkbEMbMN
Q7xEz5Mdidjzk1jpchP4ugbjjGva4LnXOpSFaenUgTAvnORdkWSwAJGGZblv1Hx3COBTzahCUYpR
ioeZRdmVJx7jJXi4YRMpxmThKRUun4+PHGBgdHtC7XUbtly96mX7fdg1RRADTyRiuXq2ofbyt8/i
OYmOjfP67QjEBUA5om5amAcvJRsZkCxgBF/pYbAIgQwe35mG82QjRVst9Nzefu9aa8KLSUZeBx7H
2vKALqO+lfcw2ORZSHSCQ5EaNqfP1GJOM0afOYC5bhDeaig1HWiSydiEAfJW4kLIFDNJfC8A+406
CRv4DM0tQ1RuELLDZ++Qi8eyekuVpnC7WSUxMzx/LroG/itYgLwL/w7M6s4qcQXdn5yvifl9F/qm
9p9BlMl0EnQCv/i1IB/7GRRYxLW3y7goNLxCISOOB4pqDVFKi7AeyYoilrdCq+THH/QMK04XWcq4
ScMFtEYON5flkbFBJW9dS3uE5dLsKxFC394p7hFORYd3VSwx4EM82zCNL0cakTOdZISSUq9uuky0
lXthnPilVKGd7BXc1AiVrrPqB43jVqLWoiiwoNlq5n7npZ8mJC7O5tjEkRx9z3bVqV2YUDT3laPx
FI2qbQLCfYCW0rfj4SIt41tLEjSopQQC98jQ+7tjN4VIUV1WfkviWJhjM4KQ0z6ArpXGNr43ZNE7
fRwBFm0aPHz1wDbhuTh05bV1QDuMvOO2yQnPnux+F3zl1i1tyUWYbHGHOenU1d8qDmlby2Mvxosa
tc2kwApQCCMZxdN1Qu4saKCwhoBcN7tTySq2V7mB91yccB7ZEp0skv9DZbZkS83Syjxx9pyqez15
atmwdbB54Ux25m6BMCYkq+kcKt3B6uSh91ZAOjWHj7KOeYErPUVoShNg14AJa16sbmd2I1UvHQgL
jdxTCZFDAAsqPvynOfZLfPGtIfk1GRM3jT2gbDjIUV9AbkG1b4vDB579JupurX0wYPCBGiq7Jg9s
8D1V44ATLIbFa5raJ/iYdkf6TU9ylEhKLDvflPYS7zjVzKCMx5aFyr96S5a814KbIO9yI8I58K7G
rBGcYAK5p/VbeuOfBvbw6ZYWpntxelT/P2WOHpyp3pqzH5nXn7bK1Bw/yOlX+WlAAHyu0jVM4NHY
R+FcV/r7nKZX0cUQubHhNxhmltLwc3CjVL9VX9KygeNtccnyKHi3hZ76RTwhaGVJ9z5MeH8gUMbj
hOa52E+6DUYphcFbHciLQGlwe+ZCq3Ep/mVrWBn4Vp03zVK7YBjE5DARdhFDa5U0OkR26XUcf8fw
+47HYn6TwOxH0NCDYArmeD+Ob9gn6hncEyX4tTJvKn/BFnj1xgUvgN4jkUT0mm6m/EX32kxwswAk
jYJBhEusqX6nfra6tzw6FG/KPYzFTKDuFYMuESzTXG20SpinMh1vxDU/ipfP5gsREVnv6fA+MZv2
vbs6Ti87TnXmBkFfLKz05/0p7saT08DP7S7pYrlpqyRjkNCBfOS0r2tIODOa9vC8lr+frezWcLcD
odAvRJpViZ0A16TnBglX8w2TfgYNTS8hY9kUvClfsdvl/BxIubdJQifiAd4BEErgAX0NPCuUOOwK
K/8R6r1/P8L0WDb/WIAvlY+TPLO3FnH6QLj5ossASrK93NU8s1WqlrW8hBxa+k7cDFPs29Wqf4Iw
/ftkUqutYKCV6O7PAblozSYNU2rYFkBjb8Ke4EZodb1kpYeO/s5TyFCTKT+TQbzrmdKdT3NvvhGS
NwG4sRcprpzRZw5U+QqGY/bWwWvutKFyinf/+08ZJIqC5N/Ol+OpiGlTw5QmDnmoc39P6GsZ188w
wIfK2jM2hCMwvvXXPXwiJ+LqI5mNqDoRq7lvoF63tcgMgJzxK2Onqq5z8D8t7dt1nvktXf357aR2
itnJbKG9p8T5wkdhXRdVnyz/QiL6/Aq1Vafv9RiM+pEiCMEelpVa1RkT/isMpgBYgiLicGiRYHED
i1VZ2y++tZKt4s57xRY4Lc5KsKUJs3J87/ii+rij/ei2Q206bXw5VZs0MjZjpx7ffFVRtltEtswL
wNxUQ8NZzrcjNFS2D4dVEWjuzDF0BpkLog8H2uPpub2clXjc+1xIB4jlKF/045K2qz/LoW3DssA7
GfVRHoYQ4aHWwp+DLabe/xIdcZapytsQWzv0USq+QP7OWcOM0X9JP8ZB+WELKSz66UvN+oGPJWe9
l1wme+wvnNgOhdQKEVFfDEOuu2ksUg722fiG+IWL2XdWJqYWLwNU1RUFsjQa3x6iqwx4BFZRT8Vp
dCmCX8cLiFIG3cd/IeS6GxI/KqF/oEQK7i1Wh7in8AhPzt2meHXDKhO3ZKgXjU9G23V3vQlDNLwj
Wcfp04Wi5g500uYh0Twt81HXaMf13DzJ5sCSUUtUrfl17lQ/66DgDP2AZp550L9xcku5puf7O6qc
vyFh0v6KrZDJcMmgtyOcUjdcWmLAmYphCK1uKqag6lluv08fyFLdkJi6le9ouAbZQ+XkN9wGWSz1
BqsDOrzE8Q024E3Uo3ijtiRYDytD2SuaYYvIxpUdNrqn2G/SM8WpA42RjPnhnYBxH6HWGevclidL
4J4Pjw+Ai3JgoaQMOxF/wZMLTh/LkOb6uT2Ui0cBbQ1hRatGafKVcvW2jxFOwCwjQDWNmNu3xyhi
eszbGO2rlHKsiX1kQZURjlLO9b1IgQf6O3+pAE2RsQ52jZXB62+1APtWx9TV7MCN4RKagtNtfgfU
CJ5EshL3DSOzRtLawb44bsxUiYTzWGO/Ec2VGtApyNykaZYaHAB90VAWJIvhT9MfGONdazbB8kyy
AdCA9jpbumXZqMncFh4mwVCRb1DA9OV8+nSr/Fn3G6gZ6sI6ojHJ5BARr66T7yiKQUAYYaxlfDJt
17n80Rs68yzIOesAjTkdhJA9pigVrcWq+LmpFtouKT5ZbjC9JpJrUi0J2ooeRpzFIjlRJpC0o/7N
wT9i12+VL07GiZZNdSOgkvLCPqvtJnkPVAXHC9jui0qRJXT8ESAa6v9lBmUaezZ1T+7+H937c+6/
fhf20x6UdySFsOVdYOifrg94voJUyxZMq/HCzU04iuLEWE6Qo6D6IdlIxe4685Lm295pI3ZfBchx
TEP+NwkQXlQHu0CssbWHxyOuAy0bjDoDfa+Qx8yNvvPgzRt9ypMbNzi6qfRB3p/VcoCgXJYXvoLU
k2qpMk6ubXkfmOj4c3153cZ+Cr08eZkIj561YwhS25CVcUjltxZjhc3oeN9FhQYTm+X+WcDXU9Ea
KmSK2i16QGDf/4bIzhWI4cgmEZJgXG+AkRDJztNeRRMZgJZ/QnJ1bNPVsLdfREsrSFC7DXQ2sKeQ
YrNoD+fICEP8ufS7JOCs+JESL8JKXnTUjyC17ov3tgDACDtRIkGmOxrCZx9I6RbzQs9yguxuVP2h
eKtw3Z+4de3n7n/BqWrjIJIdQsKIiTxeCAsBAJfeMFHyaquTOAeD4FLRW13Ko05cH76G1LyCwQVC
jJEiGjOA19uhjqa7y7MEiZcrXs1jKDCP506KLHbDFuRSTVAxOlOdVybFxeKonmLkRzCALo+nRJLR
usHp9eFjjUn+APAlw+FMReFvCH8Gff3nyZ/cQe1GHgL+px9v0CuPJ+mCSh+JmPWaSC6zyIA6W3WL
Zf+k4FemxX6iEaHeO/T1p+XSgBu4vZJxQ0x/M5tM539cQnin6OKYtkk8+iviOT3aysRmRP93uEof
L5EGL72AJh7i1M60sMzQswemyuHpRNhL/+HMARTAjEQ1MramMaQ6C3EDLFlCa4YnSZPa8xZwh1pT
1qeyzXAWfkQZxzSsHA8xtkJSLD/5BI/nuookq3UaLLyzGYnA1RGw3SrfQrkMjmM6mhCZtILyRlzi
g2dMOuMqlAIpSKcSigRuS7vJLWOOjvFP0CgRE8zNQoLvNYdP/RfYAjdV70zI8im2ph6RytUw/x+J
sBmp6JH953AkbP+TskaxCCajbEB68qzqgJ2fcYZefcdpHoc+UTNo34wo6wWtZXyQiOtFq0mmmJiV
P5hwZ7PPq/MPJXjmMalOGG8H0aC1dT1Fh7niycnelgqzEy3M9vnWBhjsQqN1/vVy47vPJe5o+UKd
INnTk/hf3lifk4VEk+qc2okybWc3ihrlD5JbbkYmVBoOOYSrRsAnRb7xxqhbaPeZpzwy2gsstmkB
H168oRcMBaGdFmVdvHtoyq1u/OHgYr5wWoZQNdZdXI4kCtYryvH1CR2gdCUC0ZQcE2gvCSqpSO3D
Ur8ph3mGGc3PZZShsj+hJxT8X+K/GoN17qjagYQkz2B+FCd5DYOEaCB2sJO0UdvtV2tP8e83u8C1
YPaP5HVy/TJg2+FeUrXTbc8K3X0cy+HNsfdNovUgUkQ1uzCy3C4VsfFv1r6dNYqszweX7n7qNdDB
UsSQH2oZ5EpREDEblPJG45BlStCQ/SSAyvSjGrd5d3yCaiGdTja6KH5OLuq8gHXTMNoCqRkxpSLl
qWgZCyVsuj6aePALU4gnhP+al6QnAPoFRbeZQD37YwrB+o37rHRYDCHlz4bjxuXqYNV+uyXbjQkC
I3Bl5lYt6UA3YWRtnEaa5xnTL62j2usAeS7ZZToba/9/YTTt8jIte3d2DFOJy76fn2eXH3GkcNrn
ZaFa6F6dIOPZCP1XJMD5uuWrNMkyig4bx2rHLf1p/u51tPBOca6JzEGBRmCw9iWLDxyCvS+YTGon
+U+z1WcMwiLXAdQEh1AxXgWL2zDeNxYgEWuQChsMAVrLm9jnWDP9DVXCbvBxqdq/ay93JM1FsKUc
asnIKVD5aUwgwQxc8qGLfcYvwbuwF17IrFi8+jBJsXwF5z6U515feEkmlnZrBdqODl3NqhJ2q4d2
vECM+SkHDwHYXZRA4CeYakUutCaH9z3zNba6+CbeegkQqNJWIfjhCfZAB7mU9Iv6KAzhE0ctqqnv
8Q3qFYWb/flptmBTh56qBrykkM3nwHC5njI4tTsE49w0DzttohgjffAviCuEPEz4OZVxdaBnXjar
KwXH+q0xn4kDT1DeRqWQZoFhX3Ruz/McrcGdrg2/xMqnyTt4rduPYMcWa4yFimLDWQe0rZXxfJhY
0ofoJc7LgruSBE1TbxD+GrjZ120qBhRtu6QmlUBKlV4GQ3IGzYBnnribsfaGkxGNmaGIbVqjO4ct
9evvQgZ2AI3eJdz4xe30KO3BNJTab1hdwn1J/Rm/1NTGmNyAUa1ZfgRNYU2+OY3ryg0+HF31HGNB
u0hmJhLtc2mcsatxSg+0oUnXIaDE3u0cvoGn/bcRMxNOg853WKFbZkyi9rgCU3eiRo1GfzOIP2d5
D8AHo1PfASwDl0M0Z3weJdccOIfsJ2j99q9NYPF/FSBUKknKIAQR4mka6gk+FeqIkqy7pZTDpnNy
VY6UN6zwOYSFDe71ayQ9w4HGqMrOV0yAQRn4oVP/gDvcA5ObPyv2r91Sa1j9M+6knVDw+PpGzCUO
0QRQlNp4Xm8CEs5fs6sd/NzEBtgLTIolOqnKaV5Qaq2F+iPGLreZQLUI2yam62ZOKL1OBCsnUwla
Mui2574DBsEqsPAa4hEApWzxEecFgGo341cP7VxkOeOPioBnh3T6WdB93q6MxJbLXAKNFX/+ysqQ
HVRBTFJjOVLq6Uu2i03PgTHb7HAF3EL3n4gxtfmENtpF4nz9IjB3rXK0snjRFH+CzpXKpRattOfO
E8ZpRPyEpXtfvgpeJtdH396qaopRgTaTyKLEB2YPiPjCCV1sNWaPk1whOdhBPIS6NRvQeDaiMEQD
2q11tEQaPZAxCZv8GlbhlSjPgD4mLRcYwssL+8hIWrrnFdaLBjX6OrzqfDdbmxd5u8GW7rmHa6cZ
s7CfSsxKUaWxPt2hHcrPwaaRlOmdLj7LjT12VwnlhjXjY5dpmgO6NSc7al/uq3bxc/IrDHK7R938
rJcDe9YVdEhIfvBtz3uGO63vrrvbVEHdp+drRaMwx3K1Hb9YopLjc2XxKNb0581tl+7dYILnAKCh
1MdF6x1EN9wG3OSl3nGQz8HmZSuBZPC1zRcF7YjeMdN/CBA8ztjGEnY7U0ragYm4dd48J6th37bR
R6QjHQWl5U+2ZY47DG3B+4DHXl7yMfr1fDJ388Ve8vjdoeoqo0GeP5b0vtqlLYyoVAjWKsP1uMcj
+ykOVEheEBBHYn6LpbZbc/gCnsM4s2sYygInzsHppoAlD4qudeorMhh4LiuyEVNXLpNPM+Ktmjex
Vzg/Hj4dTN+FKugDMBdS6Xp60ed8/REpp//9tawvwc0FJ71X9HxrwIxiq4GA0mrRLa5Qa4fsXOQu
T3SLwLViUgXSk+JxVWBSG+00sKqlKgcFUn3g4EhQA+GJWhz+TH0X495FyFW525/U8K5fAagHwnyC
h2PQumMXoUH9gsN7WbTKoc2GX9nfhCWX0kjQcyrgmz5sxqEBPVRQkPFmZJCnehoBqM2wIxJikR1L
Ig5A6lLw44CKqAkK6tmGaZmTFAsFxuXOorZFEP9rS3UFVJYF5mJ2FcltPNV6PEfzd+HRZi1kgLke
G430KBe3q0v3UMl9gl+VxtCM9e/DAWxGZwFDZptIPrtr6w/i9liSeNkTD1wUMQmkLEu8YDMQFDqD
u2v28N5Uz151WZ13ANAJm2HQjMnfw/j74URFK0XB8LvsJdVpRBPXttYPVHhAxw4si15hqjB2Qzri
g+nE/9jeY0n2nX6+C9hjv55rFcqz/mPjplitMIlvJaS31Ed/R/X9rYdAEKQlivPn1eCR37hiq2fc
yYpRcK9mS4F/LxRBTVuoWYhswtW0b79fKmWRBU4ivkgi0fXdZTqEQrzqr8N2X6n0Wg36jcqGhgPi
cROnAFwe3nfYjBVOxQ6EPLIKwmdUujZX9xlKG0darAZXUA8YA/XdvdUwp3BSVCpWZwx/V/pdN9bO
aIAxd3tI6usvUk7HuVxq5QtGLUiQihWZWPRRaWZ+8G6bhlS4Fym47Jg1zgNY6cGYT7xekEaHDqXX
DGyA8bfebNju77tdH3uF5ok334qSFb5H1mtpVr9lbO+7j1bJI0KHDAei1GUPNhY4w69DX3uY4cvW
wD95ry8tzGQ45pBJFLp1h24VcGrNWZf+Stj1bqK/G4uVp+XnLSOND2tAYjdPoA/Zk0uCoa/HwDqy
UTnlSstibd0rG7VjB5B0UMmyL1A5N6zbD7599rHnPYRemAWCaOL2ju71BDI/YscvAyot3/2V2gEs
8ggqZzTYP3esJu1EplcQaC0vZ/wlhhUZGOWjLE06BXYc8PophWpYUQV6czqkD+excSyUGJEEkk/q
HtpzmsG+HlqVdY5plBLIr0fsRNtzPWOf1rg4cj/XSYxBf1/sReUU5hZ33XHu8n3swh5pFFnzzjww
Cg8RKt/h5DJn1z1fQ/Rov5iz0yJtUzBmusW+7qIkMaC5OY4OltauRJ72/5KX6Aq4CYFA8bJcvKSV
g4r5qLDfkcRICkXM8AYjejwVgXBpWZ+dVtzRBT+mbEUgT46LrxrEHA0DxhKGfqZNTEzUnkaPEHGT
mcqvqJm/Ss3xh2C2/ha5idMPho5R81xV+t08LHCSaNFVNT/Iqobuje3G1nAdXDIj/7lHVnnEN3/p
igvkcaD9+QdbBIWOLbRGL9ibJtmu7QTA9UkZLi2A3DhJ2odOlMWjwQOD5r0HQHMgNI088TEx41ho
t3Lg87Aut8rcGsh77KSyyVOC8m00u0N2oPajmGOnL9Q6HQ3DjWH58kN0NBGN1W8IGHbulN9+ChZC
5ZoKgS9QPzJX3R1CxtitveLlFeCrQ/75hTgjV3K8BU3Oo+MPd7G6hvrvrj/eMpR0g0dY1hfNqAYV
kB80g1wx00WY9v2Qzuvz4JKl81YUnUsfgTiMKxxi+WuJX3F2XZZm12u0Cu5tBxlUxzyTBpXd84bF
IMUGhgZzl5FnxIq3iQ84IExScBBXsDchKl1wztMeTqVTiPXoOw8sViltu4suJI58P+R278zuMgw9
UpeYGUQciSzHldmAtRUyh6GN2mHqKO5bEvp30ds/8TZf+z8GT4kD+Rid1bsZ8jXl842jsb4bVjZG
YBbLdiZLfNIoqyV7UUv70Igx+zSKEUtT9inPVwSnT1Gpw+tAh84347+CW08Zo79V4jduIr4pJ0ll
v1qe07LSn/yrCPbUPIclNb+kiDT8CMxvUdbcveuq8Crm/IuEAssp1/iPTh3ZMfhsH8Lj/fJcJTC3
MvZ7V/wMKqmw2X+8jPkQGLYyY0oUYFr9J6uqyHXM9QUfCNG626dm/fhwKPa5kKTk7xdiDKuodG52
WenfW3OAOgn3bACbyt5bQqYHLMb1VLZ71BESeEzi8+uA1FoyIIdWR2/MKcdxgdhSPtEOL+Y45TaG
HqVvajg4Oh+8Yj87Wn+6TptRDK3Ffvyo2qNq5S9V71AKkMKYw88tgJk7l7bdequ3kpbAmdSE6D+D
NZDp6vo3lZGYPEj7TDLoVJ9vUlc0s1Zvwg2g81FaotvM0YsQfpKS0U94IcbdW2LIX9u74l+cuXUQ
oRQ7yHHl/uj4YdkSQ07DDxTVbCrdnqcuVOcy9LOPJwABIbVcHwlfnrrrX4brHvnHC3MaSyv8w83l
m6O7kLyoIEa8HCMAlvUSmakA02RDyPsuTjs3Aa/NZARRdMebUqQ92HpbPfFcaq3Y8k2b8S6drgse
NZayqmUxV8QhQReQ8ivWLrYDKmJdeHZYhzUVDxDXg7jj1mxoF79gqiAsJAqhfurvnzzq6QpI6EWa
lr1m6/vWTnmmmfnmM6IqX9jsqB2BPx+P+rUz+CEyHIFQa9S3loSV9omC2TDqM99RnM4U9LQQ4YXj
LhW2Us0clXCT4XTOh1KMexsg03anQC2/suht6xOLZmOC82Mxo6GUT+RzGXy9n0SBBmz3vWlLGxTN
sKAyhZ3Qszxx4M348VP3WANEv/BOpkB4pAA0FxDcr2pF5MKPDhfkGbCd8H9PB+H4TrqvcU28AxXv
Vn+OaroFEK8Ic8C+uf5BqLNtOgqZwKLmozJXqcEcb09MgJdfOqBZqPOG5cKhZELNu655G/XtcEjI
zvbG/LLL+XpEQOp+0mg8qpdiXkJDmm5SLlgbxRGesju3FtOvumnid03nqf16zOMVGjk/aMSmfrHb
aDSpElCtH1SnPhrh3DGhM3Wtksg+m2JdqwHIm85q983krS2AFrlpMpp4O3QRVPRTLX02zkE+TFdV
3vEb2eFRqaXqi6g97Ruf7CTRHrMhB6QrpLCe9xQRLQW4QaCPvgFyBf4WW5Ga/FUoIrix2+EbLCy1
mypRH3nCTg4ERt+js0FQ5cyLsVxRyroL5nFU0bbOtAtbl2wAABhGXKncKb+83zSXJESyxIrgPYn5
V7XxP17Tfr6QpTl0TS30Tgu+7aYbnk3WUxxgcgbGtDDQh1uIxanH961aYOqZ4Tl9Y/F0wxBhmcul
ZTWpeuCoELycPC8EjOvZujDyTjnqzJvuO7jfcxJ2VQHXB7qRpp6cNGfwIt6O1owK3QGwtkwp1vjL
DhgwRgqc/6QgTVus4JHv5KUaNCy3Aw0jZG9w/1C48DrIaGDEMcmRc4h4hAIfbhtbHKt6jTNr4IF5
ZaBYq6oggJShRIUVTebXDL+Qck6NDPzFQgAb0Pgrcg/GulVf1NKYhJjnZOPpmSLjrJfCeFQnZA6O
jAgJNYsp2kBpKBSRlwmk7dzTwIL982GFtsX3s20ffHAqJLCZv3rm+sa9yTXTcf/V3Atp1HsBsT0T
EjkA7ooWq0HttQo4JjGoKf8XnTGXcdOZbujEXN1Xt12DxnTEZHxJwSQy/lO51rKLUNQ5sFIA/M6q
zE++QMBqSjVWtCwYwe0B0c8/tlu4DOPfX/sWAfulVOq5rssEr68uTPSkTU5gdUaJve+6U+DhG+RM
sm5m6PhZuPSHyT6Zbx40DzHpG3Lv3bMt30sOBXHMoOjI8TkryDzhdez4wMUb02cE4NxLqieU/8Oe
4Bf7Z9fi8w6jEmr1xkjXmwSYL79ehzjbRE7IutmhszJgPgaJRRkGnSnH28Tdr56Zm9jrJZIHN8nN
WSViI3T6xJh5Gqb28+6UJ2/Jrzm8VmCotAP2TcW8ZeT/wx2W0upg+S7huC7fE8AjcwT5zQyTj1we
oCSM7nIgmCzFXwJWfYeP2DJyEoydHzT6J9v5UEW9tv2CLEf5IPeplecyXI57BOfQncbkzm/oGKv4
/8J+ft1V9e4wD82VmElnj7DPjp8tGY5sPDKdcQdUPNxpOmxcmOmIUb6+LSKwxcP6l/tl3jAcJI5C
J78BLMHtdRjYIH3vdcbDSDfyp8dFt7Z6sBh21D9ONofz/OMy0XpLLkj67KIS8zb7/dxuYMtM9gfc
B6lheSuaMfYVdBCB7Kcs0p082fpp65CPinmPD3VJOmGjRxnnP4HxVYCfehej1xOqb7ynD5lKIDzq
86sboQPM3529DwvLX38CF5OhFxX907GLCP3T/yEFqAycEsnLfplW8uhOlE9433tj8So4Nup8yj34
EbdgTHROB6FLCONVeLsFMeg6sEIZEseGO2QSWu2KD6cynKISxKhQzGNfjD2x54wHFE7ZAUl6QkRQ
cCvjOYaQ8OQAfu3GtGEbNEnLijO0Cj7O3/sfa0dkl0998nFefL1kMYKPc8/cRs0jNSj8azTrpdBJ
q59HkSRTjuXmKqPyqo4eO/66jMHFadqY0tuUOjbK1sspbDg+pwoT0PJPFvuXZBu+fkQYaL1qfNUh
fxDvCAvu/k3fgQ1ySTdNMgGPnftIHv4kUZtws7IleSRN4+10cvh06faMtqLMNicTTYmvQvkwhRL+
f9sra8CxkLjAnTqyTCcgQJ5jc2zMXFDv25EStDDFNfv75lRNdQ9FVvoKqVk282ovJG+Ojph3lZZ8
QEoo4hGXzhcptA2Y9ib29jiMUh5jzfchayrvspsmL0dHm6AipYfYxNU+0UvK2kpgZjQD7+awP06d
76D7qLnAZ8RLqQKltTzBsm30ed0Xp7ShtiYHfy+Jqj/tBlwkGm8MSpS+pd3xdOpVMqSr+u3s3Aub
jAks0PyStsvfBQw/BWRRQIA4bB7VTtKBeiokcvsYvWWJxSAGuC8S/91ORrOBgY2VuhPDCA4UF3KV
iz2gvAVV5eJLeFDKgsothubI9dYkcSRqCOlFdLETpLhODIJ6po2Rge7A243uYwwBci8yoTGJFsDe
3QmPyWNpnHED3JR22WwdENcNIbfwRAAMZTOCh6p0pFW2SQAOkUjAQ7P69MH71JQNZD1mWT/jpUSc
Sgy1khAlsgJhR1W7VbYPI46X+Dcv5NjbyS44Y31t1nDKtQ1Q2mH9IGt+WKurC3wfDkDN2UVuzc6P
EnUL2oNfp2JasRcrQ6dXSFQkMFwVQbrMEu4SMqmoXEdBnkke75/A09LJAfJuCtRf1R04kBo00hAC
zRjt3pUL39FQGuBrEnzr2lD5ZrOvN4dWg97bo/pY2+ziemV2nVcrv+IycrKgq5t8IQhP9mtINaNi
/abHJ252eIvwuz8tQ6GnbTVna+EO1f+ZO5HT5b0e7QJ/Me1g0IXzplFpFtmHyDlSHUoJbKHl0p57
9J2onJYZcxXy1xjl0JB8GRU9PI+jeQ7MK012LPajzroU7DaJNi2hhkPnc0QCprnlncX6Hep3WXaA
bB3mQ1u//Z9/g7ZDJGV6/WQMBFNm44RLbBmYrnL/HS4k8sqConuxNdJYyrihnwA/hU9Ht+ZRlQRQ
fIq1qIQs+ue/lFf8CsQUVbQUjHCobrIxMoGTq/cvtOBCW2TtOGx4pKgzTnN83MHJYg2uM6uy1Exy
XmaaBt7w/xMoQ9RD/7ESs+4N75+x9+N7snSvEbCL6mjTJGIvdeVw8ti75Ztm8UARkD93oyjSP9Di
MdcyHjWzEBS98uCGcmIk12hjkqDXWl8vRtqsV8GDs56CybfeFoKq0GbnnKeR57q/oDF70JA7S7WO
uLDieT8a8zSJa7gen6OYT1XQxgURqVUKBnl4zD8xToOcy4f/I8XJhW5tf2MQIiAVMPu+o8q5j6hL
J5bPe4kZphYi3KFJSmLZy+zWwrxQ5uyjasbz/S3tK90PYfvNYYfZMaBIKwALwwS8zlJfWz+c2Ipj
e6PsTOfBvS0vqfYSvPsJR9pReo2yMzHIIi+lbWR+HTGUZW4WAMSIJunWq06k1pJflhlfZlgji3ZG
Z9+hO4XgkluPGIAqfIRHC2W3f2dOaWAJZb+xnO07uY/Hoi8x7WC/iV1tfYv5T9TIaj23vYkRVF1n
ZVPpeD7PZwt1bURZ0UmwlH8S3Q0z7J1cx+v9Lf5VgejIiYvnp0VM+bMjeAm+c/x1ymdXPOqz5m23
Y9ijBxhD92A3gl4sM61/kFw9hjP8OaaDs28D3ZWGfeH/iI0nIyjSuh1SuUMReBEiMVszPz4Bm0Rm
HKMOsmyVf04iz9nihq8inUfH692QMH16OcZWB5HwP51Kgr+JXo+Vs3jM3IJJ1KrfE9g4wXRxuKFq
rxbgXt/xO5FoxgL27/tXa+j4jfJUsV9pWeUu/beKOS1RsGbAP6MKcxJDxwXQBO+bBYP4se49+4p2
s1wFsyyZ7xNu4FA2U6jhHeKEvCEX3I6l7YKB3taazuRkPorNmGf+PXXw77YMazpqr0zSdUKHKqW3
Su5YR/o04AnM5JUTBTnfCNdLK7WZErl63CDclehJ5WxprvxkWrjGbJf3pU7IELMfvpOHVADnmlj1
yChXhsCzXLtG3Xnd58ADXDfFztr/6uuivtgB1kAjsAC6ZNJLtSEcGXhXOZl6vRBDk/svu5QPemlZ
fnFx4pS4gG3pv/KIqTI45eqhaJ8GbqrmjfqwQqk1gQS9Jh0grAnrgxtxpihOm/8a87mNaA5UiYR3
keTZzmM/D/H7fBbSs9YWs1wBu9QzwHP2MEOFxb2DL3hXoUgnE7gwcBSup0ej4/cN2d5hSUeSQb7K
CBKZk4X4G4KsKeDRPWHxD1CIcNyEx8HApe3AGKvVYcCybD5TR/l/oZ/425/jr8BKSI4xR2Lpy2IR
BXJRyotyVDAjLo0ws8LgdwyA6L0tK6PdoxEswL0UYEpn07j7V055tP6n23Emm+Ih6MxRzBHVedrz
TOnCAzhFEWsoqLeY1GtwJWmk8OJtg1FNvVtJBRfmmvH+y7oxtbwy6Ll6rby6lv1s5rB2rjd/UScP
/RSq2ATNJpI9F+Bh0qkRVSCBcP5CWtlkoRcICKnHxSbK0U26ZAb8sxCIl6ucsLo5tgnAUQ2/C53r
o/2yOd1r89mJq2v6WBK13Ztu9Guva8234BT2sxk96yjPDKXe20Kk0/pCbRBBnczVCJgPOJGdAs8c
blEAtrClcDoQKt7xii7rSy76ninwh/RZEsw3scNYAvaxVwkc59IL81dONCatMuOnC6mcWhuFPZ97
QOfW/CfjKk6E+GNG3BRS9zFK+N7Fftd432PVi0xclE9K6LjU9cotJ87oKuPBUcJ0mN3A4JdCEIC+
flytchZUmcqfLu3A5aOX4d8+9We98f8UFqlTOgx4ScLhvAqX6RRKXn8EbXJgc4zR5RDiOnrAaigm
g2dtHVHLRE+WUC0DrNqjreUAquOEtUxx8WYRPldZNzmfaVIQEVpXha5ZfZxM8pZDWAaoLGiNDSZD
hRlu716sIdImQ8gRTKIMBQbWZ5ATmW6870sx4JJ6QMqr8whAhsfPPrtlQjtWNHQXsUseCWAu7S9z
x9BaTFHbZmfiIO/A9Iiyl5vh3vr0/Fznu/fnUT4N/KHOm3DlL4IJEW98+z1tsMfsMPw9fkjLeBpl
25FFRdLQ736JbvOVm/llKuuBgHrO965JjgT6wF8KPNN4LqrsK3e+NZtJtWqoZQk/WVOmr3Cor3uV
BfswF+hP21ZfxCAA7EMRlNSk4q2uMN76Jo+V35L6a1MjUElAq9buYXluCbUrynxT4Cbj08D78Jmr
tgLHFbgAGSYWaBvVwvIF5gNSmqkKJTkJY3Zb05uMA6EjKuB45Eh/0ISRjO8rD5KW1fG1/I+nhUJ0
7gll3ETt6QPYx9Rbl/uniqmXqWZCju5WzbM8Y5Pz200Rii0jh6knZUpoA8ckyOYv2jFOk53urIbr
f3A/vGHasPAbb1K18Mk6RpvE0q9hAerL57cGebZWhMzGSyxOeqvY9tIVxWRgzKyIkmqlZi/TudrH
orAcl5OZ+HPyQGWum8Q6/UtLXvk24Q7yz6n46PnjqqDSUN7ybGM3L2nd0fC7kL8Y9F+PahFmC4fR
+2155EvBxObQnz0jOTm2aj2CPYQr7Z5VyJokhYZpBFUVn71p1VzMzTM4ukjOGfpWFXIVMz9+aIIm
3JWdCaJ83v4wnoYTdJvfLFh9yJnbGbuHZaOTq3OJIaqNFrYwczXiBoC6MkIzdMfufPL8n06Z/kmN
D48FPKoimdSW/a4Rw8LDXgPbM8pImpk60s8u7P6ED1U1/co4CwFzlIfD26351tHeWbQZATBgp+4C
a1sUlNg1ZrZtMeD9P4PHSaoWePRp0mMHj1/AoszfkWyyo7+LMWY0hYXZO9AjNE7uhJ6txG/ftYlY
xrt7TTXGaBSNTkZoZayYp6DladwrH6OheQOQkc+ERNy1DnmkSS+w2sphOkFSgb3RY8SdfAzCAM7a
r1QAwGftZ6TSQ0cwiXHzjFcN1t388DeExaflU7/reeVHVdBD0KBZ50bg9MzyoqfK8/Z7Ddn9zX0F
SOLcUdlB0qFCCxVHmUnH4UwwQVRNNqG5Jvf09lnOuJOdTeyeFBWqOTGSQ6yl/rCzpcFUWDjyqQ4Y
coFdz2WH3v2NISK+IsSPtq8f2jDXk4jQOysYkzRTq1fFq7T80ORz7hmjwwtMDz55htHviebUY5AI
VN8ph2ShbhiHLQ1gRl4+jDi4ShFfWf+AofdSN74Lg/XP0EEFiaG5xNdMygmqbT9Po4dsjp9tnvql
Mz+QQpIgNj40RpZBVKPDZP9vfFXndDIjjkfF27IZVBsYI1ut1sbU+p625BVoiVy3qI6+NNPDqb1S
o7xY5MwIjXMKFc9673KwKGwJWFUtfdEq7laqWl3/PUAkZkq9s1TtL5Z0qKaXHHEYgJ+WvkT24iei
TYRyTtiECyUwiZxm6DpyMcUOcA/uBl0lSTiGPVPC7BE51zm/S1g/2mwMcaXuqLFocIoQH1UX1qKj
0RkJNo7Z5zp+Rd9Z06wrOOvHtUvP1MVqGOnMNE1O/ST1/kPe9yDL3Ow5u3iR3Ru6TelLFQIvaBX8
Ebx1RCbdET/12RrysGbJRxPwm2c/0HROJMbRnuwDNN0TErdtnVMK9PNCnziNY+pS56NqSJyxOuCP
WCrnRkUXEDj+JohaBpbfVTZFtIKgqUMUVL8Wu5H1X6qJFOOU8ru0etdtn0MYNMmnhpwomQ0nDv2l
CFj7K1/y4B8wxNCBDRy4GWriC8BYacWN24xDgJB6SqEpyJY3/O+eaMBwF/NpWFS8vyNk/zaZdw8v
iboHDAyURpAOYxLg2f5vmPZEUaTRi4nupQrIJI6pQx+YkjGYNfuqJJ8/77vcPhZEJPmkQZfImpp3
RiKcj66dytXLBI7vAr4hl0ruD+d6f5XDQpZbliNSSvP/r5ZPEBe9x5sV0du1HtFi1xEjvidEBFOA
+GJjRBybEqLrXJ/U/geE3Ct5/yxBK2NLoi4+7xu7SWCB/WgSIqjbgdxrVQ7SqGY5+P3h0SZVib0u
3t02Y6wQMLioMVKIBOs3iWNgPQ2zfnPCvNCXJ9ZWvEDw+loAxXyweh9CAiyAJx9BpN5CbSm6zDHo
c7RKffQugvWxLer/MGwZPpEbx3/V492oqdv7MzW670SlPjPGnGUWwpOUZHOdTpayp/MR0tbQ9jnS
88eHR7a8OjU6T1DPAyKc4WuxeIkuTyIbLzNSYyqyjqeifcdKabP+/tH5zGhDd85WKMFVVb16RFJQ
gMPTq6VTjj9NAIqKxCj2rcBdeIg4IByG2rpACge6amPHBJCLg7whcQa2ApjzfwORYipQC78drzEO
g6jlmhaeM0mU1V1mXAze8Ub6yGi2N5cUzt6AZ514iBNeFbpXChErGMWH/6scYZ4cXy9rPh8HAdQP
oVrT2+/OSQegpRILsLvkTRqUTdma0ARTvPyySvqgZ08EqUcNL/KQbNQaP2DU+h/zmiwJWvhoRfbp
sSd4y8LcxqADxYvOUn9l5ysdYgYzwDxqOT7zjQ6B4rzj57NJ7gkcp+JR4DjDgXynbWBsWzdEKEX1
lKtJ5ieoM5Tm0/FL8UCDVqYXXUvcnK/43I3Z9W3TZQ7cVXgBys5YF18UOoitprRGF6LSmun9nwn1
+rEfa5aoCxmGIllWKGD0AridHixVwWmkbhYKc9/vKj8vz2SMs1SHNEdAcDqU7b8ZnXxOwT5L9tIA
LpS9Myqydho6wTkc+R7L6NQBGUiBxdvnSNGZkM/KxigA+7MO421fZr0H7ezG/RlAtuUX6CSWK4nK
OzANwyyMb3/+0Ayy3ZIatBzhPM5tra45NUXjRlJ0QfFRLRhFo3qx/WQ9qLAoPJJetN4z0Ra4Gz1M
58ETF7DD0zrWWh7T50AtekXQNTb5MzzubUfWmwNETBReK2xENdGthxKpuDYB0o9BuQoi/JGcLjs9
DmwJKMOzUive1LweaF3ICHnYO/bQgl0rGqv127um/qutcVSwuSilIodpBfOOtgCjPFaEDTwxYBD3
6Tg0fegH4v+K1lcao+C6Wr1ozlLZsVBn5yD+DyMrdLB4Fb+jHhi0pFFD/vGm6JHps/JSDwzxWym/
2sHYaCI3l9cI1HXrnsiXo2vDaFacJOh93lqrXlFiQoLHq22W+IN+kp9C3uLueZFsht3V+HOaPTjg
0NoSmJeanQuLrL730OTBr1aOEBTRnacnYpwZT0D5ERNeCLEpoAYLeCEMIQND7dbAiE3r5nR6jVkB
phB5W89/7LStJyfDgrAR5fs1xm5QK0f2ETkuASO2+KB6VfVjVyv5HNqL7BX+J0IOM8Xtk9vn3IDu
ZAhA5amSbmWMmQDmlQdY7kEo7JjO01ciEh9kuHwKcWHKL93QT+GD4UBAzZwv2RobpeOqSi5yUXt7
tmUHZg2Z25MVLLCWwYTV74+C96FrgOQIHtI55sktvACoEjjtf31hvRLVC/iNPJclYzLb3vh372+0
g9h1BP8NudbsrPNDSX20fE8Oy2Mr2yzh829RzSri6swPYwhPhj+IeQ7OybrM4RCfDTGXq6dJ8nVD
JtJHOYzIhkjUmtgEO2nBPNWkYzjlKgye6BC7IMUTxSey7Da5r6l5e35Jvh6VoErf/HeGxX2XVn9z
ey0V3gGCTDrFjdZNYXQxrROaQPjPEqkq15QN42QnV8BNicBaqzX5FoyPA+In4FYnrmhVxZibLLsW
jzNe5QB7MFYLXHfJjBlsDsTtbxTHpM48o+PhOCw9jGltBXKPmO9+XABzDJ8UA7bwJG+BuYvgZ9t+
vVYNI0ZTxx4cs9IoychT/fSLpTiSx3aagqIbty/l0Xa+njqoPXbNs6dZnJwGBpTuwYh2N0hbjNmS
uVMWylHWoP5jLDMJ6G47orFUSLuw/BL4+OPbcCNf7wLbfvy3KAe2ib3r1bWDrSk9Tl5E8WobthXz
W2Im+TClZmdloqhZE100jb2FI9d+fqPytpMJ/lsst0f8PyLRKEI+xhdT6kvwFTa1EmgOMeC8fMJD
N9nXn5zH7IjxMnVEaZ6Cuqg9Rq8wXgbSNwy+Bb/qRXLCjaPAkDpQHAw3TfhKLfsokuRaeeqPbFnv
Ia6kPqqrCcfNcr9hlQIH38qlajwitbRn83WLdra1j13zlpYG34XAWz8TIRlMsmoXUOmqIF3hx69t
7WUSVkWqEmwIUFC7f2VqBBUsVAL4sKrXHYi1vPBCvku6QGsv9NxpHriJoE0HjLnEfIcBhv4bVQs9
Cc7GdN0z472i4M6YbdTciOQL/jipfP1wfTjWDI+ZEhCTgYu6DU8Etc7siCTkfyKLvMk8xGr5Kjbo
xSFyx0TtCOTSkT9sZUZEU0/iuBiR8R80VJVT9AJWU9n9mKqNeQq6L6x/Pke/bJg1XhUBduRp9np0
UElKaym9ecAXJQO2PNOU+voXp4E/yNC5Gt6JS6jumEdGVACTaYaH1+rJyr6XzUl+5E88DNqX30FF
pbPoEK9bMhYiaMdK5iy5g8vLQtUBq0RxLI1EzMhYdDZzh/DjmMHtkthaUjNP779bj9/q/hn26NMf
/pzSr+Ofago6LYnPwfyvmNiwFmezK6E4zVbHC3ns137ywIsglUrAC8LA/jrOt+ib0mWi62SVphZ3
n+OaoV0ZoiA7RhW/it2wtwkzSqwmfrorOyo/vbfOFsGMwJsYsIqSikYKvM4nlXZq+6I86J1yaWIl
u0Puls7vpLDlqlcZs3mDcDU/QNALadq8lHSH0u9MV0EpsTUQ7ARGP6HHoln9ep7ZQcGZ+VmqeUYm
/65gpuqNaQGIC97+Lcla/u1xCCQiCC4Y5833amz8NgM/900YL2coZJDOb4I41y/9SL7bdh3ozO/M
v3sXJ0QOchCgHnIJ5wctwxfK5hSH4TlMyIVnaMMawvAk5zUb1VCZK/Bkt0uXYthC2WNLbsT2oO8k
0qhQf/WKggRH2nQQJAGJUctteoqk0AOxMZK8yu434GKFIyZ8bbnS8hXqZ5pbsSyvJiTm/0K/sL57
tdznvUVuV604jZHtcx34uv9gSMGXcU5bW3q7mTa7vsQf145FoggPi86W6rCT3jVI+Vbzo0OiQjBb
rwYnhxGsfG2U/1M1sp0n84mjai95H2Ngqjg1fjVQbdKK3iKUERjG/MeTY3dlkdyCzESIKDPCXdWc
plhb84qlRSmSHQp/nXBHsc7zkNlFmhzW0cq+cQ3tQIAqdLYea6BmojMtq+he+obOkVYUhK6/o2uZ
/gglrnJ+YE6QvTo/27tsx3JC0XRfffDxNcxI6KP5drSzaHVlPXG4e4zCO4x+PzmRomdMzqfr9REq
JTnTGS0u0Igk3tkt27MnjyUQ+N8cqcFUTkD+YN509ju0a2n5YaC4JTvcWXJIDAwY8Hp/QTOZWssO
GK51Anu53ZteFBqTbPb7ii3ShcLtF5ysPD28rrpbIt4uoLmcxmxy0P61fs5e1YvMqx9AQqK9tAku
O027SYbuJLWP9EfJw6/5c6hEREn2dWmtVBJlqseYZzxQYGtRvovX9yWO1iqOxJjw7lzDMyWLrCv3
wjT9V3shCw3xepvwQzgefha2sMoLw5HvgnkpHD0R+nm6HzyxDfgn6TzwRNEvjqfVS+IdkH1zMTrk
BJ1O6+zWr8+BHHARQohkzp42eaSgSA7Y9s3CPvh3mPEW6xdA/PXJP5U9d2PJNVrRfLd/k8y0RDBf
mTjPdfOwSTfJDrgSByrwQrYHC/1ZlZiNWRUjO4m4pZKzF4mGqkr0EO/ZlpRgECj2+N1rwO9IVjSF
2EG4hEdkPpTCgqfV5AwN7aIXj8b3nWqyY92w8Mb9gcXVxsWmyCgvEZZjtGYpnJucCNOzWalOnzxf
Ze9MAb8CcpwS/dgqolBbww9YbJzaAbz1J7N7IIUQvGiwDHpOzwkTs14KzcohNqs2W/aN0NCVp+aZ
yDsZdBo0eUkIhv/nH4XGbcFOY6qrQ5lggfs0jODT5INQ0RADZku/EZVNaArfyRm/9m0Gl+Ne3cFH
n+qCRaTJv00BBLh7MEd2nHxlE8sDG38VnFMRDoHIAtNKSv5Jrwv5nn7nBQCEsFv1pubE2qZKumAc
9oEa7XbCttQw5kZcqAi6oU4UnGw/DpbTyn1J8jBbBdjdD9dai7p0/k/27TkCVmEhgnfZCgQtxfph
PYwDrpPZcTBZuEJ/ykMg+Ig5LwD2YlZrsKw0rsBN3rL9md4Gufr+DwNqHPk/ixy+kKmnI7LrfC/L
yqeY56JAgcMAYtcHm9dm5u/IOw9UiU+9WUUKIIstZFlHIuTFkUlZVCd2cuq+BYVE6YKpI7x9c0/9
R8HGi1HXRFAC3Su9TpWi0fxliGAvFQWxX+0uhCD5i/Ja6LGNpI+YKLBmlPuYEHyXupdDAW/s7yzJ
Rjcx7z/ophslZHlwg3Lg5jHOI4Urm9rtTBMlMer2pbpJob2i/ubCadSFT/twIq7S9sQ5ZkOrWWVN
OcG+NNLouKKK/XMwZ/9bX1xVmRswnMLy1Ipd1UKqkwbTDnjyUeG8hMyYQ46lshd2JwSMHdr+L9je
54PLeKId7f1o+BO7W63l0KzGcpfRj/UjmeZYaJwdkrxzlTfVvrUQSNem3zaFi5CaM+MAP9IH92mu
JnLtNzGhs2m7Kk7wtORtuwZJmNlLRUs8iw9daT3Pv5ijUSBQJOtovMnKBwaKhJSfnxFiyOkPDSnW
UUw2YYDTRdNvga96xPo+Yjuq2qgVHfamb9ED4czg7o1YfFaF2w2+qvqgwP0BXLj2GIan+voSSSKg
pm05Rywl+Ps6k6rf5XgqBrUisFblT6y2eh2/EO/P/Piz5pBepCi0KQq9Hv/MCY88VPyM6P4y1lB+
eERtkAqQ4YRMDnaQuD39bhu5iQxH0nrzDws5MzBU2U2c8oNiHvJz8ZZue5UxyKvgTBSN/Mq7V6P7
A+FnM2h+LCAciGThq9/XKFtn5fxsMtdT55jrhN7Q6kfP32NJNy71leK2FvccKPG0p4NR3QgALuLL
TA8jKejIFbddlh4OJqSc00FKNmWJtxt+MDOSb/KEvfDJrfazz1hg40gy2UdOlLOoW2tvleVUPDYP
zDZmVuU2qsewSF7rDmHSDKNz7oxnQbu9TrjOfCOdKpZlKAtJx6t3Q8MdNWVvHqjFJFC9ki/A8ElN
/gT+zVzJs17+NBQx5b4KyV8hnjPDS6JmY34Jlb8d/afMgCMeubUCc9NSETLu6oKkNlsylBS2ftrY
FTr7OwSxQw4Okxahy3Lt7mkKn6pjMWCLirCrVbPWtms/+BTMlAvvR+LDBlQMaN1zkbOIEW8Ax3uD
Ayo+xS436+Iho0itdpJtkcblPZaQk72619pDkR6g3M+eKoHCk2QflzX+4jDefeSV0sJIVmksLiKq
lNly6H7BXgYUkq+4DQK6c/4twHu5GLcpTJJhEyAHcUHe2SZZo4Mg2+L+nJU3I1lMwFdckWQMKcv5
rxZiWBuy1Z3Csyt2iTcnjBBTbsG8keELCQGX9ljAOk01psvh4RNnzvN8AmMzVuseBquajG3IYN3y
99Yardg3JVI1oYEjS0P2G3aps8inwAQWjT70TtU6HQcdcSNXH3x7QNmgmZiosPV1iA958wl1LPjB
YUer6jg+ONicVD8XAqZstvgLN2HnrGFAnqp+ISyxUaJcYWqLQ7fBL8Kq9sIfEwGVc4or79N63P6i
b4XN/HzY01qg+7JokAqzG+aRU0Ai0m8qBTdyzb6FyZRVVZGCmbVhcWX7qXODBenYcdGBaMg0mWeq
lJTW8s2gxIz3UsXhygmYWj7F4tZjI02vCuVgyUiCU6L1BOMkLD3zOHKFO+SugNydRIHjDDmFgG2Y
DPpOj4wrFKqS2oDAgnLRpGdnEU/usP5jLp8v10RR/PfdGs1cGAwqeVNrPrMJ2u1YDgag4F/A39Pn
zXGdUCnQp9GNi5I48EGz6Pm//Ifw0gnY6VYu+cIBJRNpT2tTwi/OOPMgYxakeKKjtq70Pnl95WMA
o5Ro8VJcC5t0P2UQBi59H2wByNDr4217obDo5ld9YOzDH8iHJYuI6LaBUUkOD5ZmJz8rkYQljTAA
tSQseoY88bgYNGYWFp+/0n22g3AO0JJeGmV7I3EThYJy1Q9MEzuRfeOgjCW1PnMZsBmR6M84Nys8
wbZVaoHzrb0hpPWxf6ZJE0bUd6ROjgyiu84sYE4rKqGqceVfnb/miFUVcSaQ5FYjA+T/4nl1d8sq
0rM0ZPE4J61t1N4/EMxyDnSOym96gX9xWjC0DnrvoDR8qO+zLKseVN5XuY2t5ul+wxrfOGzAgGB+
U84B+KZdOtE/BAN2BvVnWTdPPnazHgz1DJWYthHEGYzprNuHg35kie/AO6pizYxHsdl271nlvhAo
Vfl2wO2hYnxvrd67hc6zjPIoN7vIgIIDWXY4eeEn2g/P58HRxRHA20oNoQY1GSY99/milcOuJpsV
RNNRbz01ipYu0kOEDVQFdEzGp8nTEVL6XHko7+YbOeiAprqTUIMTYSWlSgnbA/L8f2uom0NDWIM4
eO9gkO3+faE6kuuHFC3h583rcglp7rHGCNJIZWqOXaHvqZwCTuDN9dhmno+hqtDUF+IKW9pF6A9Y
2wrnIaf/u1cKQ25dr3Eme1Snk1lFjdfO2PKlmDKkB0GzMk0fK9WygD3chQI8GnrIQLWH+AyUco2P
ROMchRBbMCI5BkVKNmvp5vyhiXuX6BfoTnRCGe30dCaIm6dLqwZ5Xib11rHkWXruYMI+dbYvMdqP
IsYjOstQ8K7G4j9OFMEVi/XCIv+3eQJiXNM+9kpORArbJAakt972rB3oy1i+WH0PQB14zRowrE9F
gKGCbgxq2pjvR3RwT+pt0/3VSzQ8m3GL2021pXO1ipp50FCcjjZVG4NFq87p11BVRyVBP+aa1Tsh
nZaz7DgA8X/ZFvXhVNPnbwAREvfdL4vJlSqDieg5QzMJUiT105pf+9CDN8Hwa1xIUC1CuUhZ6FMj
cjXJ3lNTVNYmyZieAqu1OZvOK+HkiS1VZSdDwUYMiaWOMATaqaiK2nMfbz6RIcpi4CEnhZd/WX8G
A3MQwZ9MrdZYHifUNGCSnjokOTlkb7Mc2SW+c3lkyPiAQ6rK5KgmcS6v1IOEOLWDUCJ3MTjXyqnr
HHV1tnaXzZRdQ+ZZvu2HdJLlRhlzPJ+cZom7FJL38XdcbqcidWyQkMtsAjRQU9cvqLQA8Q+XsZ0o
fk+q7JmUybESXyJMRRXOnIdP8OyRVD4+PHsuFnfGIaGNkLeVhxqPMhyxuiCfwf2mliD34SxecPvp
QpsagwI5gbz9OQohiBL5ZhOZAvlDjk0kYjvGXlFTrajnkAImTIH4y9M/lDDYxE7VyQ2FO3Yos6J+
cN4aWwR/NV1wQgjnxLAl413QLgn6+/8oTbCOWcHPJABym0ocsp64e+I2p8cylhXRe6qcDEDKC9LC
87M9EHdrrBlQJrkru4LMemr9xItufXyaPWCe9pw9C9uGI8v8iK9lnRZUYM/Tshccx00CX3xuC+Tc
FgJSnXlzpi0qqRyQQNnTdX1fGaQIRZoZYu4AyX4NGypaSNtFYbu/l/+89pKyZC0tf+/ZGYAfMkoD
AEOi3mQ2NMNXEyEraTJq/wZZqbvIQBNzjRSQMlFERHHB2+JfxWFzbDu5i++mhjyWCVeTZQNcO39G
UfbByhZ1/GtuZ508Dx1Yx0iaEzL9L4vJ/unxfKq5/jphZi7wrcas9sv7i9sUIPTUlq223MBVvaOt
R0VHHi+byQF2PWkswzrI20n3+y/JzPfQy6Gk5F9TFzOyLypxPUyyszGBo+0IICwnhDVZqPazDyfo
GTveSWliZ4JIyP+E+y9r1eq0QZaxVvkfM0xrGwEOcndTvxypS2l0naJifbnyTPF+e+J88fRCFqNr
oUIQ2sAfgmQ837T7G4N3unwWYg7fH3NGxTnKO2vyHN15L5EM8jDCuT1l/TBUgfT6EVucAJd340+T
PUs6Rp4whD5Uzx8eFP2GaNdVVwMz286IbZ3CPRxhvfh58Hh7ni2p3PY83XJHkqNDY4iSf1IsW7JJ
lA/nZKrDg/BWK3li8T1Wj6SVkwBczosWWjCErf/HYx55DdoAre2yNyhNi9HHq+XiWdmpC2dNO85q
h1pADsNMnlsJ9Z2vAJkrIutwjC3pfi0C3S1M4hPk5y1g6s4K4AKGUe7bp7j625+PtmSErQjtbvRN
Aslg4Wxkuv1zKkQ+zk3oQgAqj3V+UgZWF8UGWsD9Fthz8p7c7sNj/zNZebcxVONUp+SNM8+eiUBf
czmdXJFMWPw6E6vtjZQbkr5ZAoCygQSqmuMlExD89NTqfQiE47qM3iWQqYFZMpiS2Cgbjt31cFeR
MHntSEWMFbXMJEibYpWl87SV42w75ZBBmgwIm63ahafogh1sskdvy/yt5DcwJ55EEaVavgD3jhyG
X0Gbob0Wt1dg/gQDftnOaITOFmX0uIA9/qv3HzEFNvPtHcpvIe83Jvc9U9NyBEzWkgAOPKBdK7jJ
b6dfSAvj9Gtb6pjolOcu6KcQx1e0Pew+Vwzmq2KwDHtoNaHcRhaRnGX6zntVZa1G1a+01y7AxKWX
5XH7PE6UNhCyNC8+OO/ESfWOr2aGRfUgp6Ks+D/3NkfgRcw+YAKFG9ez9Ozs5eP6cWswuvGfT03Q
JBQay8xU3MWXogWD+B2pp4cRMwUSdjE/52V589ENE7cnbDn7KjbLYfXS3NkbmaDbRj8oQPJBq0gx
sqIl+OmSgmZ3xy81kPQ5Xj3o7oObK1b7TU3MwS9Y/bNxCwq5t5eqOoNdnY5AgdBgPtd7st1/EZAW
2zfHX8OWQjYTNXPPmYX6etZUKGsyz++CyESgmcdcfda12zb9WqnpBsZnlC4QCtobRxxxiiGVWU3a
23yhFcwjaxmZ8l990diJRg95rQ3cZeafCib4QsEnidar5zHqtnMsyd6DE9JnpbxIsTwAtFYZtoQn
m1Z5JaHaEzmu2y87/d1fx6QGVw5sYbw12TcSJ9wgNqRnBdOGsgNoSa5mP+OZ8CO2Ho/R+KMTBuZX
pHH2f1cogLZi8YJUO0mgleP7rthIzKK8NaDDQ4mBRptKq4k2PgcpsunXpSAIw7eFIT5xcZmJ2PU6
Q5rIMvt39b7cQ7Hs/6KI124k1xFYpoNZZ5XufTlbUvWqcgIsUVG/LqdD5x0ygG+NXWDFW6PDo/Sf
N/oVK1oG54w8ScUYxhKX7HhQwRPcsB8OXKtwiPmNmViEkH0ORwqx7jpUrGTVqbYPoZq8MemPv2zE
AqZxagC/AYKEkFwZjH/yD8tmAvPB8DC43S+i0oUnKl8h5iLzfoGpjBXAOWDDebDgHDQ8MMa8Nfik
o1SKXAyDSCdrqUrYZWcnRzC6ea7TXDINjbJJByR1FFNt80AggVvwWYC2js9a4dvipFtZo9V1ICKP
eXtd/WPHmMs6D4oYSZX6QJ4U6t8zhjECp+qlLnYnp9l6jgiPikiE7hwnc2+1eOchNjTZts3MuO+S
DTJYHeH8xIZ9SbbjxvBys9KaWDHvQe1vlXOXdKS6RloaRfYfIG8R2HhCOxNiAcAhjs7sfBb2T9J7
LkqrKIps1Up56GbEMVY3dFg1NRR0h8mYWBNV+mEm/SobrOSv4rmsuJRZuE3ZUaRq3UUCy5AZ5MHB
rSaw2+nUAet7QtHU0bT5A00iUoBTN59v5lyjs2Jn2+qxp2vSB+J5bUNnViL9Nq8uUTCUPqpfDjlx
zf8iU/p3a3fTOf+kojLReQy93i2jfXq2MNITvxWEmi9mvpwheIuUsA3KiIgo+ucmRkCenTfoUKG4
lpD8iZrM58poVON5dpvQJfddpCxAcuBkl3eTtzm0LnXUWHVw4mn/hsebeD7laGtJ64TNMLHrt+/E
Yrhkq7o2jRdTcwksVilt6O4gyvVgbFx+sA4oh75DM3tpoudDtKQ5xKhB5jx9y7DIN9p5Oev1jyDs
Gi1n/4Gj7hRtdwO1h+9Y8p8qghsDhuffNdKscIx2Eq0EFkBOv15Lv8cIpbwgAbycv1thRicDNbGS
NeoOj1Kqo5mIF+rpg+TK28bG18a09B/EIMm6+aw5e6vH5HPnbBuP/ADsziwHh3tFo+0i1VpThMHS
oshkwmvVcr7JE3HIOosunyzU2MOM9wPxJLGpEnUthbji11aJRwibzE0nUlSUO1irma/p2er5rVBW
+6k4tyM08GjUe85i39GrE3fCxFyi9Jlw0R7i5CODbVc291ajWL2cN6lZmOepIjcEGCNsAFDA7n1M
MEBbjH20W0ue221+ZIWg3x1soDlyWrQ+G4udmKZTnVrm00E5JnfaNKjGRKJeqWz5t+EuldrYp/nr
esl2bYbPkzFMxWu2HrwrRIq4vWRhQ49wv3UyUAamYWigSpM/vZHJrZNXLmD/ORHTNqnvZxlbK4Ae
WzsGkaZglAY7KSPZUYJO9pCqAdOXahxpxnIfczTM0EwJxbz7T5k6djgJ+mBPPZ22Lyrh5Ya/wQvl
FuUZc10SjuXJ1oOrxJi+OeEZs3NV1GYRhTzIV60aDFooORJ7dG89k7czOPNyEBWjdrwr0y6N8nmz
hU30YoTopf4Y3bYj4uDe3dRU/FfayRMEKpVcTiCaVshud7DlOHaH8fALJO4dKtn4sg7oB8LSWDWR
ksKyWEyWtagVJZmozAyIymqv9JxQptWJugoYZM7hjMtT3wMikD3e2OSyOPDGaF1Afkl7KUBDyeBc
vgx5cEJf1uvzLVlqMjuS0VX2KPtIkt1NoQh4adcRDER5gcNCmvkISL9Cv5w3oHKiMVQ6EGrcintT
ZOQYazHJuEcpvDBB8flMHwY2DB8ZKs9y/R334UYPLt8GQA3QjJIxFm3Yl3RFJozvCwywjhH7o2Ia
b9SmRbMXQUPbtwLj6ci16Gz9DLXnAig4Zw08e0VPYrt/buA7bVmL+wJJ8khjbDWns2ZZ8fZRiPPZ
3c/B6wh544yMsNRQp933sallXhBb/lNB44Myiuu9rk2ADE9NqZUrWriRWY9dq0H2DVtmak37QcZV
OTgmJsMdfHRSV2JhvT3woz/hYHZtrweHucsUe65AQNH0l9b1lvGLcTUJeUVJ7DMMCQRocFp35ujz
xigaFgrIj3J/LL9KYI5CEJNxWlwN5Dd04SsUQoFNcR/ex1Fhg09RwObf/ByXfoWX0uKo/u8kHzv7
i18Q45EhyPhUQvKh9MV52kwOOI4yInaMwcw9eSSwo8lzhOy7Auj8PNrvixitvQ6dCL8zpuHYQ8WZ
UmCLZbsuRPUCIqsz0EpyLY29rDPiMm7Z/2yMD+mFWjwVnRTxea0HFFwgAVp5mRY9bztJFxTstTWy
/z9FXowpX6nv/srPvAuPOne/LYOQXdox7J9OCQp/75/VQ5u9izfjRMyy3cTmwoEca3Sv503JaEg0
mUz1W6vhb4ymBWY+WGzKd3kIYREzGxRIRt+XZ/OHLHBCg5SBNMxPx2Vcx6uNwTAoXjwxpgQLBEvl
yvocf4EYXJLHZqfHZ/EsX1L0+MutpUBXVf+/WYEA7OEF2oeqlRmQ96sUqftpeQoXlyCx5PFPThjT
ckMam9Uhu+rSmkvKNL8iyUBXHISi1bjOvFkWp1CZxC2YPa6Qq2zT+CSrlETFNT5SzMBlrxtgT16F
cpTMwLiOO9BIHICnzklYNPlZIlGHbPuMhU8Y5WiRldo/jdStALU2fmEpLp2Tq2xo6hRahBOEzMzt
WBiHsKLG7H+85kk9Z3MbuuYnWtExTC9wnTmk24x+sa5Z4/dY0MRD4GqYhWOnupt36SLyXTZFg/qW
g52ARf+z6dqrYdrHntpEeFRuZDGmWSEaUW/jcVdDk90eriAJoYIzY8oMnZvYznDhanXkpvLWlSM6
T+Wy44nGljBsAALjnaaHO9i/Wj4GlEs4OeCFwZ48241hmyI3YxswYAIfjePxaSaC7I0/log2asPX
WwyqJmumvU2xEb3Nn+Rr+qR7qkA2L53h7Vg1w/z6EPjB8/hGc6+ydlknlDpAFTWXF2kGNHLHwnTO
S2YzMLnFjmZmSiaNV2oQs4QUgzXHCEug3uXUWD0wayEMydAFBVvIfrI/kYaEFISfpHPhnRk0P+Oz
L6preqBnLf6k1+CA65W9VRoKNT6IpRKW/yyfXd+XxVcCCUKv0c8L9BSmx1EKMK1X3/4diY6xs6jl
03EDd3awgLNsOGnPuSSXO2NzF9pfJ3aHloCsUDahyY3flA2Oic5y8+QaMJrLAbLFWcgKaq6f7bZp
QzXskFf2p20S10wBKhwUDxwFm/laJbexIHNClkTXHNsMXrRTZQVgRJNp6gVnIn1kcvDcbZkbzH1z
2q5F8QsDxkeeyVmCz1zp5HunXfadPDjphAdb1HP4T8CUdSBXzwNdBWiquvLprLHli1KCnK5GXE3k
AZz64GTZQymt83TseWuBQPsf5tTvI9Fh1MMZKYug5PVs0uUwFU56VzKpZxNYUp4pbSHqS+7pa6yQ
EBmyrv6jLzC7Nwx61fYQKkMAxX4/eIYI1jYVro+f+2S6M/tmTE9bjJIzhSpJdhukrHkHV2CcXXWu
QJvr+kc6jDCTojUwccGZ+VFK4NQhI04bei9XULa3gYnKiVfRCe/awMy5LFSDIpqfqb3WojVDbmZD
8+b2qZvn1afuCpT+sGTRf2zSjTAJpqmDINfEBWgpiIWHXoxKTZFpZdQ1pz9InrUYb/qqU/NIrgTR
3vcjnRVBUwbE/bzXVyrTE8SVhhjlKHiUbaXpWofCX1i8YAYUFUJonMRefKHewdlFPX4mRsJF2/wu
ZphOQrzYGNOn3Us0AcYqLfXVHz25a6JizJYJDATLhda26I9pyA+6CAyPqICjx6K3ScPflYHZ3YDx
6RtsCyG2UqpGCY/KilyqPmpPoCWcVYwuHXT7LBrcZOamMFD8bCQ/mh/mpEi6ycYnVfR331gH9F5u
eilo4t5Ke8NEh/L/ubOEJjMuiTC/Pt9YyJ708gK4Yi7SnNCmE0RaOizPPW3sG2c2mMgwCisQj3ob
UvjAvlIXPLK0h91G+mp9YdV4dRN2OYdz9bTN7e4ESsBSaCVHZwfhoUF8TKQVuu37Ef3PeMahHpQZ
jfCTkkPd79WRuUn3K8L484kF460N+y/HTvwQuxIzZ2IaxxkNGY2hyMv93dpGi/ld0zk/GW4IbmKS
EeQLobPAxXgAIy2HLy+sKbz6t0GLX5lji6g3IOHWyznyk+xbo1cjHKiQ7E2937uLPqV2tM4abz4k
esHX+Q9uUBXO6C+o4muBPkuoNQ49ViB6SRxeQ5sK+/3gw8Tepj4iwcmXDbDKg3WUyzhggAL4GY90
c+rg5I1ycNXSe9FPUKkPpSBQJurM9eAPgeCdveLb5kSzzNCUEXmXqXs48FU5WShmU2VYsSc4kvSt
EGt/2jpCmVRLURjlunNPpPOkM3eYUeD7Ac2Z9Kx2baUcOfe0G42UEkgBfP09r4LWy0IXMRb3oqHC
Zjf8ItfeZm2tVrga8OGgEFav28Mw1PB3tesZh0O6284yFEgosBkiSAFO6YaJzwXozL7W+WfNBn+0
OvKOPBfnwYL9k/jXVGw3WQ5bjOWy1MU2fdiHWKxrCEr1bqrXytJatb92vCfH96DFFSoZn0JdaFBW
DBjg7f3zXkRQZFuGevUkUAOOC0Npwy/UAHrrZA9mIAquOTKcXneGeocuDg8kYA9bGZpLXkHIyc7h
YpePqAvP+GnqhBwcDor5d6GqGc5uDPd1XhQyVX85F6jPgilGqIRwHrHto/JAPGFyNzw/vcwO0A7l
xW8Da6o+irUCuvbpXwEELpCfQP4X4460UeCe8c+at3NE6PW2LKdP6zcFMVPjE1mywA9yxOxx3ZJ0
k5FUqEhIdJcoCpEsZqDg/nAnn5EJ72EUtSgY7DmFRHz3lEC0Sb31RBM/UQ14wa6qM5h+rUBZbJ/1
lp10kg7wJfL4o+5Ff21O4O6hdRwL0OEtoglEtGd0SOLEF948IjXhHN6mQ/cNJiKeZMVcvKZgXryZ
8hb0+EU/GDamJaVGDqmAbSQxbbMu7J3KdILhIsbXW63hiHsa8Se71IXIpIGguykeEKN4VU3Jxzwc
ygc1jtXB9y8GkvCwyGV4tyGqUpjeyhB++7huHEwjQuevncqSWg/vaFDb9eAY2Q2Gwk0hj86kwqFm
Im3C1yjhkCoMJTa6C8R38XD8m98u9Cvpv+Jr+ls4WdKUk1BPoj1r3PQFmzZvkOomcbXTgjyBQdzA
mYH91C2+ncrJOetGWYiyxcVQ3TGScezGA+30kD+G0e1myG2kqvv/vYVY7WLma46Ve9x44upF66WJ
C/PtnNERjIu8Es7E7x4XR8+YH/uvFNGSBn86ZWTSijk2ROdj1/0eGs6pMndkWu0qmuZAccAsFhM+
yomcsnUhH3zCZjCMl0QoTQfLHzWGmqlLDdlRVMfvPDvoV5kio8ARH78f3YgnSV5OzMZ5gE/e+bU3
LsQ/oM1fyLybeQmQlTosRGXup6u+cfhM/QVyZwryDSSoiqCC1aJb2+kClinyPw680BGfniZEGtGT
EgneVGMf1uXDdx8O1wi7aPM4XDn4YsDMnZqPhevGkRguka+YMFVNX2W9jOLMSkpfyVnnegxScP6r
mjG3ppjsjjs1lAle9lm/pE8mTnTp/lTpEwuI3FBSbktBAxQ7yzkPpTFNJdKFoqOebde/9v6uQmEi
+/bnerCWNwribkD0dFKeVyMMSAZljdVJxG5YL1z9aT8gs/mzdKk+USeycK8ET7oHtKul1sCfyDI/
3gaT1q2A4cKGWK7p1nvJvaa45VpNclHjdgemEgiXbz3TtwJtKWfr1p9vSgS0JpGyKETJp3/HYuI8
ghWLKJNB5LSjtzAgeoP8A7thjcBWU7M+UBTWk43wSpmPaybOWRLX3ClKK/zxuHwZf8z0VeNZkDke
kIkGZI4jYpHwd3sbxuISUC8vcpbM0oGnnZLdzMXoib1FxykQwRYn1t/Y8wql2Z1VMsGrWuqX2NJZ
I8sW/KFWDR/x8XH4rsrdzFsoASw5OJd2nLcOQlkozvP3LIjcUmLZNMYl+8kNf9S9lF0Q9qewQTc6
/ILxYDuiKNqaj3YEANTpd29XtizrAl2B5wIh2w2CZCYvdR/YRCqm3pid0xFr83r+GJ09+4LmyQTa
4/uy9obHr3w/G3tYhUU0FlSsTeZlCIg5PciUHN3RtlnKvEtxfCZM9NGD5JL1K/gDhefhk/AERpRf
oEjL+a+KYGEEx1LinoJDaV6w7Or/6qX6Qz+9mOqm8BU5lkBvokP5oXUIo65wyU/Hgyk3lH1pOMVn
DrbyidEdc7Hi0WADzr0tZdt6na75RfuhpqdyKRcWfFpDvy8w7ez1MW5NAyMh8Pu/NuvhYct+SOJe
/1SMyR7G8K0mSCdkX1b2wSRkJjfayJBQpxWmimw4baJqU9hjYn4JSxFaewJxL2U4+hDA/oQWPmfF
oWe28Sif/JXFyTMwcwULbbAC7EheAl/vLGCGf2giBUxzk97wNq0ZvIhovtd0btDiS7ZGSEdLT4zc
L/ZwI/uNO5BEFcgvoiJP38YpuUA2j2sl8VxqtwUdXo0I1AacPtKmiViVImzHd8VbXAAX5DfGoylR
S6cL+MUdYgG2oZnqylYq0qfTSz7lAK+04IpkB3oLqAZ89/pUOJt3lDi2nkqj0M3szVSMQ+e1NFK7
FMHHJpXPzDa2ZV8VCBI0QLwc8scEP+I+Dpf40yp1B1mTU8IMtKIcmmTrKmH71x2uMZeUQAHe5+Cy
JQg2Dsi+eN3Yx+RHWsshKTY5t7XoAdOA//bxDkfYshxHquq2j++5ttRol7UCeC5UK55s8mNKdBL9
PVqlBSx1Q1hpZoRGq2Kth0rTpHCqN8YiASCTGrikze7meWnJQz2ZdsZQasM/u0eVqSOT6GL/L5OV
qIgH3Da5yrdnOtP5pK9Vp3NQxrMAF5rA3TkUEqD1YoWfVWyPuJhNDvG/cdSXdMEzb9GVuYWRHhMF
cummmeyvFJerj001cfxRhmnP+iB3bRse7eGWvRG/9aEkxOcAJnlEi2Kel41Yo535GguI5TcqAllX
/zPxcR1XaBMzVlFn/C4ohs7aP/yUDD5PdDDBnpZJ2+f6fCPdsakHa9T/564E26FaxtLXNcycaVFQ
0DrCmOK6MSfoA5zckA6QkCVQuaAXpeymo8+W+0SX0UMro52w3HP/GLsTxujVHbCyZHQw4aMokbxu
rb4JaXJsZ3M00GbYOXCZaUPFgmAhj86NqZGaCLb224jPQT8mfCtTEOH1FjXDskkzw5bWZt+xrz3A
AmKOjhFxs+KGpt4kguYbdi+WvLiaDeWc5c6EeNBvTpRz5J3OHNpp07qrgvF0Us1sJck/npA16JRF
+i1Yx2QTdDgY2u4mT86xofSNT1//cMf9JA0Ylbe7rNkB9Y0ANtipkP+Txjg6xmi99030uGxWe4I7
OFMMOam7Pxmkb+4VuxZem8nuIEJNWUHVHFU/16BcedB+CnlcXhIQqDd9kHMD/BpQQVn3hrGqF5OW
gJ+jHe+UYihlZQRp6QLpyh+UBZ0IWRBsV1/vDQOou4kxlx4Y8zKAL4PcJxMgXB6euvQN7MzHNU5f
5tagG7UCfkqWiQKCHgl8xM4Blh53qv6vPh84xtkBrQJ3IMGv8KUfPyAMYjzFNtQMkvGwG4CuEk+a
MKn6889jjxSGpd+pxJ8haVJxvm1nJxD2FhIcp2pDEWP93FWHFc3Me5tv1PAcaRauiBIG/tKdBiZb
H92FxTynYC8XlaWhJZhRwv2IdyxEik9BHFzJyoKcLJhS45g4XHmIMIOpXbp1v261vEYVB62oEg6e
cSAkXPUiaVXDYo9hwcPyDPyMwFKZLfuMx5BHXrHGRxU16wkNStaAEM3uUQcE+1MgOehfg+m7mUnu
bu45axQ5cBZBX0Ka9ZJ9051cIw1+NA2TiN7r7EiZF/82kkBgN8M4wVzrmpRTJ2y8pIJWuKBMqQ1z
zIbxecj4AtbzuO0oVm0+CijXr0i6c/T+8zVz/pziOxhxNtThDMM4LCfgSGQng6HwVte1ESC6LNlm
qdVBD5KDLp2EOMQCxK9Taba4zTrVA6fsvCSwZKFAGIJOiSTEefTAwngs9xCIsMP0+lRep9a72Umt
QY7W8zeE+npjNA+6GzZSeDCVMFYxH/CUDnleg6tiPAsO08fY/lwa/bUFLsAEzEYfocVF7dDlt2O2
KcYsMomVLQIz6nzxHD9p2aqxCGTgr+hx29EqnH2Fret+blIdKgKKPbu8dM+J0oh0tGf1tOqnNEKD
iUzXw40266v39sHmFrl5Q6tWkSdEDMlmelT/2B0m8J2zZrDYW7GFqIuJpvGLeQq9HEfVQkhmSsqd
FMEJRe3TF+KTvr1GNPoGcCf0M2/m6mjLVZNd9Wkw45NHZ7/nSG+0Caw1QhfU0QUUHehLycVTaJ8C
S8tDh77BzlswrclM8nwhgzlSHLtjVjuCJlXQYejSmGdWTRW5mq3OmMxPTjxutCJ7MAEBhK4GDDjz
s5eTeL01rCKnoS6GmvPbzu4n+Z8YGrarUei/3+7xIm2eKlXe3NqC71GGPjbcT28UIdWRQC0czGng
yUI7z9VGwLHNPs9Ec/jUzNmS8YI4c0fLuD9tx9FXBKTP7o5yc79nQQSFpNcQvGcDn2uWcSlEmRZH
t16Bg9HeP6/wzGJTtVDBobH+4Etw/HA3MMBjxqX6pCK4wWjGiGhy6Fr/CUk0/wmpaLkiWwdIWITZ
GARE8rL/ReZrlo+9EdytbMevmzBMHqfYnPGUAUFIq4lELj8/pNQtt0XS718/4QfL9wWqvP5o2BRB
U1nukKn2p8BqIJHaanB7NbQ4ROs+BEzJ1bU51Aobh1a2SPGiKT/2Qou1zsvZKgdvTcjx/9lZx/7i
jS5pf8h1K0scmGBqvLg2zajHF9Q1E0yHGZNC7SmVt6EukEW36d4sy1idiZ8dU8ODt1wLWZjV5BNM
nOPPYCGwf6z3ACLfs2e9vlDDscWxaIMENLNJaHhEha8vEyrnTwXLeSCkEpLJiZyMwxKvIytG0pLk
wF3DQ+Znj23nwpJFxhenMlymeFL3pk4AI2sDtGmC4wVvxvZQZipUvNPpxiFOufbgAy4uOQ4qEl1J
Dy2/K3FUvH1U87ypFAXBh5eYN9cP+hgefx6b4nktf61pk+85REwayH18DCVqziNVr9HEU67iUVdr
vdueuGHPSXdpAq4C/ZbhDaS2YY3gIFlEghObg2rZYSHz0L9GGdJg/7luGetr+aXhuoBKq8/5xrzD
BqGFz9X+LPQTXDpU8oi4N8TkowfxCBtcUKXyHeyDyYZ52VL6xrIW/7Ewov2ASP7kI9hFvrwtKIFR
lbzZ4t4naZJAd2/1nzUyJyiUyZJE44OlfP8gYfiQ4501uL5mC/4gDN4O1/qWOGf9/kHV79zeS6uc
n2AT2Q7Wp0s5ahpg6ntAjYBMw10zX66Jg6HUHiHsPRlrrBi2OIOQY0nLMbsVswJvtQzpOG4kloNT
WFIslkWF8fF0BqQubcMa2eMiXAw0sbEPe4F6qKKfcBVgHsx3y1YuhSys2w2mULfM5EatvU56FRQC
6Ly3zfwqmtD7pPHFkI0u0lvFlBg0aB80yPTVXGZGygI6YnAuD/weRZ7WVhoeusflXgm+efGP8le1
uC3uA7lu0aQPa9eDERJG2lCc1UU7Tmet2uZLn7i8FVlq+qVlEf8DfDFTVz7Hfffh4gGKfRWaWC0l
GwMo4hD28+AMN/1ZSdyOyeBlO8Jq+E4f52SS4p5flsCmwnUnOR/v83/2BxROL9Cre/HD+fYwKu+u
35q6M8WQhW2EPASlHCmLLpSwMftFdC7kG1GRB3I3/C167BaSt4o5ylHDv2LNkD4h1ofjPldxtEnx
Bh4emLIrQZB3tMOzcFaBz6bOUsi6yz7U5AcS3kncr5kvkaPDZ8qZJ7rpDzU613uGfk6v3FUy7Jse
6NdZ3/cn1fNio6TNxH3LpkNfQxi3gI7TkxV88Z/jGtTjMZzbka19vtZOAt3HZSgZYydyh0w78uNN
ll3kJEaKFq75yoH47Cg14q0DF8mQ3IbUtQwGEs7R6rxSSFF49+1/bblOhw1rIoItdoXsi24gRXli
kCx6R1EJ3HalaG1FWsRNfk14Z7LwpmFjISnfUWsFDoqpRahT3Yqfd72jo7ztGWItnTHhlqrV2Znc
2XTmhz711HIKIVHIxMRjI8JGCXlw3+XS+G7ExLDkUdThnw9NPaaceJjfgXzdtenV32VucpwLvaYk
51Jgx9laLvWfKcjucO1nSWVHU2t6kmbBkLdEn9fRGoa/C2o7ixqK8mf4HwjX0CkST0e2u2eT4hQF
fRry1/xz9hltQUiGtvv9WjVF+TtlfiOH1LbMBx9HMI/YOqTPnMguFVXb+PfdJ88qu05kG/RL/kaw
2/KU0WBk+hNWNTsaR8V1xaPbteqyTSQxoGH86KfGi7AauXf8Cp5UNn3jvePj4vNqQ6pEjUHF+aOS
vrajl51NfKmEhXrrAdjKj2228KV5IHOIKcN0bNsCWQ/kvjgqKQ6SNX7Eku2DRMgYJky4CHwb5OjZ
9+sO6a5EiEdn26wjzcwLXc56eke1YTqLBlFsCg67HlPf7fYhsJkYU7I+YyhFghHOqEA77bF0hWEH
FEZpVTef05C+Sr9KhzAaGW0o45FZFGBn2HrUYRBsahDWkcjTCXI4sH10i0PRu7Z/q+2PMBSSqoBY
6/Dys3aO7CoH8o3STQz2M943g98wn1zqj5b6NwYIgNyBFOFzl2RidVNEAiOmBzK66QyphSIaquNm
a/nla+gCDn7KzxBF+1z/+D3a7gu/jdkbZCSr8G0BjTrzxfu6/LBSDb2TyNaCIYRzvBGjpqvuPpN0
q3co/V6cfclhk60LgonvQeLzYy+CSCzGSr/HAGoEWCbjAxuuq0axR7feLpo/+Y3gB0QCgx67aqGe
D4gpw/lqRrydzV9yk3j0dDgF1QHYioB9XA/z3m1jgU5YaFjRo18OkghYsI2DMCM6AVJ/LNqsL7kd
LWcd6omOs65ONCJea3sz+eOXlAuX9ShTr4Q2mtqjlvudzcMdPxkHkhYKV6Kgfs/5jA+Cqv8YLBJG
mW2gzjcJPuRVlmzvKxcz5lP3YYn5GJihpzTOr2tGtiwZaSKPbIqmyUTaUz9Me0see3AEtV0nBwB7
PdoXSbyk4BWxUrZW7Tn46eHTWs/P3v8xdZvhzF4N0JFN/YP5DKKvK+lO3xZwNHREp3lWnuusHrUK
+/+oNi7wochvmuj8u0BDRQaY76tLlWpwaqWKYJQck9R9OOY2aLeL846AY2UfVr8d3+SMZHOrGzZ4
ALlhm49vbbfXI/OV/O2dwdxiTkbXw5mZoSPJaJxz/SfRfOq7hxpF+7MpeKHGHUGNlYx+KFxx03bi
/sAbgkRWT/UiS70egqlHPyPR+BtNZWXReaIxOkuSn7H4ihotXWKf3bXxdMakWnPfFqcQRbK/TGwS
AzoEs0Nu/BZf8Z5AL5ksRnnymy6aYqREkYmpaKItKjrJWbdbiXSvdZtAIdzoB0Utgj9hfh17wG7i
LuWJiqWZNphmlul7heRxmCau3Tz705HdhMwDsRnq58x5s5Vugc6SBo0cfAFGRrO2n9fpRlVwAyJt
RiqIj2ycSOGXTGsEqIK+A2Bbi+TgxKBzoKMgf2wbhbfBT9Y25Tbe7fAL0dsCAJAjWsJHgKNQ0rjo
O3m4UCfvNA0Y39ODlsAEhXzAvrN60NCPoIIlze069cGNtsdG1z7n2k36wbjMtHAVbCHQixZ9GOwS
NCRvNoQyX9IZQPmz7Iy4Rt0RCGcvlogyCUijBRa+N9uFucjCv5yXHO0dV6DmvaeRjkefnrFiZd9X
Y9DQjdRRQ1aDg7QnLSCWfwGLncatCNlZKgwKQOhaIZPS61FitffWyTjXzig5yXe7G6AXlWaGPn/e
PcD6ocAcSxj01jMGE7keKv4zAXRZ5/aRgfxRSRfP+CSVfPL9FaVqS68d4+pNpqsbQavNxAPYX7u8
bRBtXiHvDVJjk5PjeeUFgza1T+wAiTtIW+Ur5SJxAO7h5rBC/JUGjZ5y4qGbCzDYG6EEGS0ulR6x
JQ82i6dWqsVesmB5C9CLqUZmBcMvHLic40JU3KYs75QjLc5zxg8spnWI+Bwgyjg5uW1s4i+n5o5A
IqkZj4WlOPzTZs5F+/2G8nMx6Th0BS6A3oGm8RNsYvBEpWYJ/mwKh45vbX8I2LS6Q1dv+BXg7gKC
8yAypoCXbxXONDQkGLDQldkoHgJ10vDHBVddbMEvFXXz0vbDS3xU+k1IzRtei8faxfLiwmoXpCel
xrbVHygTKXIDGsQsCMyjIVlybUPnPR5HRVGG3Q+GHwf7UqqjbGpoS1rTaWGuA7eBSu+YOhhVnUAj
S+44yKCRCN5+nSAK9i7qtwOFD9ynptOk9Zf6g0BlDGM2ArbM/riKAvIS/EvcPKWkrl1+zUFOJnGq
G0S88+SFnY1up/1XSEKQybsQOY6eKdX2eyArk/lheMk+JTkW/NEshFObOtpJmucVVe3gG7WYzDat
aaVqq6mc62yjteAP1tzrUi8FKeIaSHob5dlJ+kq0UF0FVWkxwA1OCYDoP8u/MB3ANJZw8hR/HWMJ
2umS/op3eXLSB2ccGe5zlhYhZSZMCYzXor5COpPlx3RqDLvkmBy+SpAMqwkWUAaTflICcDd1TPVa
NNQd6hxRgL9rOxRhOkAZk5PzwPqCrc2Jw5HYHEmlPlhSquSZbSzlkmhs3F7QtYfaprdOHLMrM+jT
b0+bSZlp9zCp423NvFfNsHrjqedmwPh1Vv6F66uAzAtxDdtZomUVILmNChNmpf6Ug3yLF09D3Tpo
qJkUVZmqjJM0dqKv/mdS+i08vIWgpi90/6BqQsnnf+k9kmt2+3fYBRtsRcV6cDQhjb2koQh7Z9FG
ztMnSL1oL20ZmI5SnkUo0oym6AVHsjPci7D5E7dtSotMRNz/AQmdwm/dJUvlC/CL6cEmK6THCwi2
9towk+OqV7vczU5i5E0G9nO9xckbEhvccL7V2mQQTJS09gTIAmp5FxdMiMYaXff8z+/iiW7vlpgs
BZsBagL3baCVh/RU0z3iw8upvO7A61EspUygd4kUaRNKzB/YC2KuaAOhchy/WDEpuSMTL7IZMR9K
YIm9wZko1FrdZ/bzUYJp21H8htW5vDUyEHGHesgKp9AaWp3XK+c0kxasZiLbnWu9igISmFlqOD57
Eok5p8XjQkxIdfgtIzWH0i7u4XD1NrF6BmTdOWuCH3OOmzjC704BGmcXD/hS2n3XhgycPui4pKR6
re6Wx67qw2H3aKWE+251uhyMosUb8mOZ5FVTQHzcpa1a1EpDD3wPxRpr22reS7kueKUdH5RED7ms
3zELVPbFAI4oH8zt6DmB1S8z6Ay8ZCrMD1TA7mmsp8Gv0Ky/H+POZOlsUd96rwbY29qoVI6qDI42
j0sXcLCW1Tp3EMx+vJqOY5Tz50zo+C8Ojk00nLojcN0G/zYTbSRPJBBpZHta/gfIgvO3DwyKiY50
k1GUZxjMaEU52FZR/r9UunhNS7I0i5tQmOIEfqYUXX/FPy5fN3HTwXQlCTZIr1vujecbJTVN9oG8
uMOVMfWsvqpcTFjLcUY/Wm/XEkG2dBNSA2WHamA45ntszCeeS5FrpCqH7cqgRHcAkB2jvMAqOeAS
S9UvsoAdoGF0GcW66Hi7Q7ROodeUindnP/OqCzi9XfCpt4+uST2+MEJhhLJ1aLjYtW7QTup8+6vf
Rq/+xoKDGT0ppq91l91OFCEFTQxuFrLUzwByze3F3suCojxv9AZx3Lg1+jcbmQcoAKsxdw4qzbFN
qjsfG+8LZ+aT/dBAjK/ivwNAfEj8C9E9G87sd1vmxKQV6NZisSuhq89n3n7jzoZleyO3MGaP51Wr
8PYR6lVvWpxV2eo0+ZUDM/2mu3IjeOHaJDlOWuR0TPeZSVuQBJRurdPcRQdbtJHcQwZ0r8et9MLu
vKWY9K5ljpSpnwHQrm96lXVQux4E8zTOBoN3IMyypVUuaHQ4YEhrivrsaRTVxzGALQ/pee4IrGat
gAYb9V1ZlRSdF3NpXO7JHpWPfIc+ko4EST1M586l62N8ng7m1zXvhwOa/xvbO8XFSy0+d8VuL8JM
rPTx7X/U7vnwv7a6K8n4aJnhxXvqHHeUmKWTIoDt7QxZtHcE4qPRn9KzbUN1JyZbU1xzTvlNhdaZ
Dbb2ncg5USeEUe2KCPPRohA6ICwrD2CaUP9IKoujbmkev9O5G9GGF/ducwScX+STwJ7ARYJLnsT9
Cz06A49k6xHZKnhhtsBeZh1iqd8nZk5ogMyr76PMtaNpq26+sFtbGrgJRaSMps20MQbuaxIw0A9t
oCNJFXCQVDnsBtgwQOs73Z+XeSlHJKR5JokHl26peGVvUlMpCuKkD05HbBKG3lP8WDL0Li2h4tyv
nlab/ODuEpqSVW9p0bV6RmCIjXFm1QaGhyVPJxHISFgChdFaokrJ/HYSDWorRQrhZBZVBtakpWEj
gGJwuuOLPMog6NZ8P+Gd3kAZw89C6COvSaJBBN4az+sA2Shfk5Yze8rf2DaXAiBfe/4pWDD84/Kb
/cUpMm+eLIkDvL3PvHoFAztZOFveXFUoRpsoSBsblxJUNtzMwRgAhd0F7Ofb7Yp0DRc0522G0W/L
hHZkbspVG0bHq0c4guXw0zBL7YXyxP1IW12w47GI0ya+Zcu6s9Swi0/MDRNFzYS5502MdMGYDUnQ
1ba7QLbI8BaXKPZPiQD9LsZgEiGWa8grcsXd8gSZdmYeNIUbKyXBJQ/QlUT0YCEH/oWsiThtb7+8
JNI4D6k07add/ftT9tuRY+y7kCyR6rU/OsOJcEkuvt2AQkwspgZ0xWy6aMXNjrA39yBH4A69VEIj
nbiJnmpEDxRMKGfMpeQK2tEz+J+sMtbVYe7Rs7YBKhcC+AEOvBiSxLDfJbxz6h/uclFQ5RqewXbR
154qJZbZBqs5jHxe+IDAWMrhDDnG6BA/UwrBnKBAQ2k3PIFj7QZ9ATKSHPMcHnAISrjOg1EZG3Se
1rGo+x/QmoRmyXdq2J3ipv7cA1anmPiZIozdhXWKiK7pQsQjspVBfDOqvydBGAth9WPuAThRwvex
seXGrgmc9qPZCzBandYzLtnmOHleeQ7DmXY+y0+Nf7u99zTJhrsr1uhQdteRd1gYtuBiYgf1pIbZ
XwmSRig5ZAcH8SWs3LejSHpZo+9BfeSzUkjpjdudQtCN7SDjrvtXpewNJk3z4TEajzeTOHvXe/td
p04WkHjGy/1rJgLrL8qOTsTLb9mCoD556N2QNVGqhSLr/2HDbgPckHts5U60FVD84BHowAlouHmg
en78bL9ozGlcNo7tqAkstQ+vaYXGG0YYx1HNrDs0BzwdcR3Fkmm1Vxc52lH1bpBs0vyAxs64FRsg
ZVwQiq+JNM7Xy355hP1B+B1RJtxcYtRAPN92Rb8eVOJ9bUmPmfdAJn32jBRXhbykQFTajSiSivnr
4gesoUdGfOThcXqPRZ6pGIjiLzYyxUz/jbtUBkB0MVrMMhHDxhQsIM6VuMegLFlZqtnUSqMG081l
iJF3tnuuqMoUuQD+wABRJwrmJ7u3QKd+apyUGDFQU7a0oYg3Zy1JTgfxR6calD7T9IKcf4OMHXtZ
oCzoWX8da7z3RZsUy8c+GtwPU0qQabjsdf1sibhz3mMwfonuzjQc3uLIXLQwlkYEEWDo4SC/3cZI
CDvlr9sCAsswA+sx/8We9yzmi9Wd/nY93GsiS4brmJT+6Ad5DCbCral5TxLSxHVEeB6Bi3RQYQNz
NQlGCXeYtelgUiEe0rdvpEd3rLWVvSzSy1X59hM4PE5DnpUcWDykwMALWIeZdQ/pyvLiRoc9Py8O
CSyf4ddfhpDoH/6pc8ltxTpRlStI66DyrEw1nME17nWNIrt6/E+z0I5HnwffOgTRov63V9CTydYL
WWY+oDV2dPkjY17kh81NmKWB2UDMTYi0uRHCGIJQNdY++XL5L37gVN52S/c12p5YXGIx/0I12lIF
ptFWcEaNMGKuimx6hWh3iAF/c8kZvP+YCcin0H3YlUIIvS3c1Fk4uG+kzFO6avV5iRtDqdx1k5EN
KJFUtb1YPYCrTdlnYamM9HB6nCZckoCR7IEKjveoBZaRa6kIm0zsatlbYwGltCXy3AmxcHwKIMXr
F5pPzmZCacXDFMkE7kE9NaNUSVdFQ/bXvI+hIK9uzSEmyeGVsXDcB/vJ7oaS/U8SXKEPT5objmOr
X/H/oGJASNKOU+Fsdxl/2W5r31jM9gPu5bqQvQdTq9xEwoFkvVp/XFI9hE6IdYatT8cpDm+grB0K
y77TTABfjgI3Ow97ErEHLsD6ADvZRhl/exXUFHDR8JsihVA/CyGXVO+Br+CILk8TpvK7UMpzcRYx
aURE0CXzPEwJNrM/EQBIaIBsmvSRKb5tDyU1DWq5A7ap/UPFPdHNozw8CkmicUXSUh4M8vd5jOK8
8wWfoVrZ1u4z5PXkBIjS24de2aZzPR4pkq8lmIPppL7lHp6mqw/7WvYl6/soc0gFSNZsXDNx+zbi
ndhFcMcaAjOrRp5ZijwFhnJenR2RqI1H5g2dYHG+aY7IyFZ58Kdtt9I2+1NzUxwejYRZBgubrMx2
kZPP6uz44pxk3+cr3ce96FeQ8Lmggqq+OaxQxoRyq+YcVUjVDg80dcfOWnAr1H+BFA4JXcl7onzj
u5328Je8SstpSND/68TIGR0KB6Mzz7LNNrNgcPWX/xmGaqtEzttgY6PvM2PHtTBYN46hgiyPREeq
FkYQnemMxrY/4MXrzPr0a1f1E+VeMXX2Trz+oxAvUAA/xGenDhhM5xINAq1FUtWzFVevvi82a9uV
nTq+3X5oP0p6e2i1M2K4iEJ4TKQpNAOBdUoyvhIEXFjendyhksYk1F1gmb20pE/NU/kX1Fi3HtWb
5r6Sj5YgqdHk0EMxFPgKL3xiIUg3T56gAIWZVILihC/u/gD8bMjc/dRlzdK1utXWpvFO9E266GlG
bj0EhEOqpWr7DOCUAwC2RrUg8yUecq1+W0hcHd4N2Vp8O6kJu6MY/NWbZBaMOnT4vbZ+G1uuj3jM
0jL+u2fLBZ2Sx+YVUb4/UNMFVwJX6pEfMzUYumIiKePddAiH869oj3yKmCEXER7N8T4ZaTAyvZ3e
3PPlIe5ZytTdHE9dU6Blujpgbt2RVzkwRlSdXf6rn/XntyWDHRT++ExCYsXCwUUnbNNHWWlwfZf/
0fNW3opRe20azlZceJsxk9MXGA1lN6KWYLWxBMt0YUdF8O16Agzeoki7u1lepASXzyey6P7blOiN
WMuRWbpREPht2zlqk4SEyj4DnkT/Rnpy6bWjtTRd7yLdeZiz+5JGtlVKwPbPxIVED+Us0LkfYNff
+ZP8O9LonkLfgjFLAESQKVfSdm9+c4CP/Dkty6wI2zNrt33lCW6mfQbSGcI4J2psBxQAvecCqwgX
T3BV6LtKOaYN0i9E1gLCfAj8bZsNiKl2Ld/a+WPHw6tnxblkcpGLC6rrsZnQuPPRqQov8yGBFaxi
JL96ZM8tOaZa/bPFMPvJQPXEDEUBSs3HkTv9MN1RHf2yWc99QTqFGzXC/btzy8/odpgrMj8wnAgc
v5iaLD6hAFvNiId9guD2gNDA/pXzOIWCilqkU0YALW62xqWbFkwfZw1zz/xUUcYe3CRAiMscSWa/
CGoogyHJNBu25FLyZUwTvrcwowGWO+BTkl2ktReP4gX6Gb8UmSiLGY8IE7u7heauwMtDr5k2u6t3
u1kaEWzT8ULdXo1IuGFl258iOKJq1O5gve/jEWpHJ9dqC/iHjC8nJwwxVglAZWn+8yi1tflPzVFH
Wh0oTbequPb5haxtfM4yp/H+CMPyGbW22GRRAF8Cy3CYscyO5DU9KvPe9gAhzJVf4LaaqoihJ2WZ
4OCVShllFBGyzkvN4RRL0G2uFccwJWuIEpeKOP5b8ILKhmZZ/RefMGVL47O0lmRGT2clcDB7HfJj
EVjzDPUHTCOCxthBD30HUjOLzkRjPUN/L61GVcFwa8LaxUOsq/PvCLyU1PsaWV55GO16DEPYs7rl
KHDyqE/Ms1qZ3hGKEq3Cl+wi+Hvw2cGKCHJm28Hrt9jYI9HRVqD27d0VH19j6nGwzoawms0YEAXY
OJKjQNWcEmmY7YPu/QeCFnJ2vSagpCYOeMGOV2g1vhkMqYZMXo+hpYihw1x8eIj3gNm9VawEZUY/
nfINlp+Nzd42iuNN+0PcZ/zg9cQd6Ptp7oi+kAc1SaQ1WEZJmqVm7q7Jm/aB+56ARYIzsmcO9t4M
/dokY5MEtAi7c7GvH9FgF9fgHfc1N/syT4ls838k/kLwhTUKbzlf/WJ8u7iIZLoV+TomibhRnhE4
ZVVQ+xgIoT9ed03ZX4ASg69ypUAxWmR+IlZFIV0VhIvvMWf1tOu9CSP3S3bJEfCO5plXvMUGyBcw
rgeds5VzYtAwR6qZBmIzrdcyTuGaV5z5Lj/fWNe4sbV+dimLN+kPuQlH+A67YJMNZYxKZYMJsU2Q
tFDBcwVFgFpFkWH7VwVvTGKRvl0qY4tkQpcBbzkRvJHejGq0rEbsgcETh7TpdCsUXPEXi+d5nCuv
9QPLviP7q2WgTJk4f49hQoLqFPNpu/INqe/5eeugdF1ff03QZrtFQZ0MbtLzy3atBPuwgSt1Q8JD
jn5Ztzt7ArM8h0aWq5KTT4UIlZxW2XbdFvpAu1Gv6/4iXhjbMgXdh6lnqaBjFW0y12y2/9t32MiQ
vwqC1Z/oH+yoTbnSHRauMFykFIQyW7/wsMgoiwKLKgFI1hStT1kDQ4p8UGk5+GDMp8aSECLi68Av
+NOL66f3+1ljXmKjbSoC8ppvE5gF9FA6R63EcFof188P59TwEO8a+bLFADSsI3Y4C/FoArQMAveS
0pRsrqpB9vRkroeN8QwViOulqV3MNkCP/cZ5k7FyglKaSch0f63Ps3y7CWNNZ8mkNiyimyt2/swY
Jbb+4bii12Yk68yTptB4bN37Yc+4esWE+vWuPsc+Jjp9owWFRfT6Gs27y2OKZ1Td4+XszyvBR/gS
qilYfoAvLGVVO5+ItnZ7P/CG2QJ8doh3ksbEzloGLz7zuEOTk4s1Q5KDy1zAIzCr1ZSb0xwibgGP
7GXtiLjcOTe9xqiThWp16+z5fbslGRqpH4XVAhHIHGvK056U+qRVK7Njyk0NZ7lhcD6jfPr635Hp
tM4d5MYkUwNbWWSfY3qyHcT/bR1DUmypjS5HMI8DL+lX3xkfgJlnKLgTBmzWdjQmTlDKS3WUr0P8
tzHn+Z1u5nNqFIr8jJV7mTA4jY+plf0DIAC4YhT47T30Zsb5MhLAL48g/p2hMnePYlfMpyQ4xX85
ysSfmI8P05crM301bleGVcetL4aP9gWxZmf0QJ4PRRAb4GfKpoE69oKdnKAJJvOdUkfy8n6qyOun
whzpE2s2eykEnow5vk94WgrakzHwNyN5lgWNdyEbccZ7AKQ6TlSckOHqEGcftn3vYSCewR/4tatm
BH+kW99KKGwkKDnhh2THH6R6clPUxrGVf19JC+ifx+i61HH4E9RvuATpwnA5Qx3LwN+i8uugWBH5
lx8aYgzYgfHJ9Jpn6oiKRZ8p/G1FmSExQ7EAjLET20tlCgXQZSLKDvfCKxuKAfElieaCNzZo8loU
bF6BU3b2A4HtxGP8xN0SIiKmNMI6AUViQHXLxPPbPZdkBXT+N0XqU6QyCxKRgwag2rBMGDznKN3r
OpH4wHbTXm6vVpH905M3hZmy36mqQIvI5TMa8PUm251n+ZtJ6aLSAJ7iyWlCLpqSoy5f70WDLvR6
YyNuxov64gOJ/qSaYQ9kWycNS26E+35q7LWEZ7CtN43p60JHqiEWanu+Fgxb/EgAF3AAgK2qkdNX
H4648wYOGD4kJul2prmEBSv9vWJWZ7UXTSoc3qnMCGwTnTKFp4SpkoWU4yFHLRviCElJeENmQTbT
1oiRZfpx6D9Dp3mj6ZEBOZ8830baGsnfvu/9dbVshmRETM0R4ehjoPK0Vvg7p0OekqEBMven+d3G
n4Idhh7LQyyZMQ36RewmCTTNkhR3tkf7cIF+/cH9k5l66PSjpsyjN8HCtVHzT8MB2K2+gEAQdZLn
2aZXCAeFXsxf3FXcBDYy/+D1GouI062nDci2e53UkNH8Px7r42czLGkpurtUdPpXi38riG3b+9rq
U3KfqTMFkRZl65LoelKr8Qioj8uwOKtdLmTuO8a1tPjGZa94DkCNt/LolUbQUhc9bXHSHsueQN8M
cR9j/3PXLsyZte9CXD0yDtN84p7LkCpsoiNsEGN3bz3y9QmwbQJ8sUuAsP88ADrVyrOD9Ca+1Knw
DmGgoR75VA6u8r2l5dKHdioqWW2fZnQmuJPxdk/SY1+F1c8dcUbDmC9Irg3Jtcj7S8bOqh1Jxjst
TDnDsz4tk0NBRVDM9siNupY4nyyvSrGeQA2ShNU04KiYyPd9VRWy+gT/ohqRYuiwObpakzpqB48H
SaUzuzZTGtUZnrZqN6We5o7S47E9CNfcf9C7oEfJ3TdicgxTaQEqL/URDQSBVqSyWhyF8DpPsUSA
THA6Orb4NlJ9eehAYw2GqY6MnfUNpCE/C+e7B80dYbeiTs+eiACjc+AzkZxmdDiGAqtqzbN2lgvf
ZQZ4EzMOXCf8En8S027DCkiNi2gl/vJk5PXrEpbcLHNNjw5Z7luZXMo15zQXVHkt+SnoeI37EBWC
s4EEkFhDHCSchH7UTd0T77MrUIqF14zk29SrtSpctgX6a3HLjQ9Geh4OvTQaVvM1hHp0ZwEfcQHh
v5Yqzyn1u1j4xfZPIWWdM1AzP8r5PfcjhGnfoovShEsgK18GGuELcO5SkXoqTX82TAp88eaGUe6D
ygxXUhS1G0xIMQks4h4UEUGYwXmhKa+DGXoKiLozrRtRN1KzOaAs9K2DZN01lT6TjYMzikGJZmu0
dMyJBosub/yVTUb7dNbnNbxdrbElpU6KIxfqOEKwQUYqyxCczUdzeMie7DLUx/7dDJJS2oAME7Ac
DAg/yFpqn9SdDG6iKyF2rRsSnUeyz1XSl+zOCDUmg6GMxDz4FDAwMgYIHKB6ou94iPoAf7aEJXYU
AWALJupOYgFT0aW56XcrRJlqqq3Z98CCX/hjJ8JkoRLs2KSY50oGmkgsEqa55ETAhMbqGEkDZa1e
xt2cW3sTnv800q70aZeqcpOdW3q+M4sqm+r6OwbczuFh9XfmZWU5dsGujDv0CPRnihKQSWlDrUCL
pQxJMi3neNelH4t9VYgyhJSKQTDqHRJScLybjI3KJyMQ1Zol+sC/reSVE+68E8HM0j+hDkNcEnqy
YhP5EQ/M/CkQiqYI3Wb9zrYKSj+nGLp+ZdHtfSipfuNrjoLvarAREmF4zQykxQNBN6GID4jMy8Hf
qfx7ULFvI3kqizYFWlUcmNKUKfLswD8EymO4OvWyjtMxG6uKAUuTYPrgDt81lJ+vGtTSs31NHxfu
CH9i8urO5LpqzbQYCCnzXgATEYKYTeD47RS4QYyEdp7/HWXH+HknyitNf5AL1s393S/zpqiRrYSx
OKEVf63ikPnWttP9jgfHQ9c2WsYvpavOiDTh1cPhFjxaZdYhHTalmR6EewvDi7+iPxhj5S3TCpwo
dWnSAkL9z/0Nw3aBVdLwBKReIjKBV2S879peLGOHquZIe38szvL8zrPhslP4gphkiHmmvk3GGltn
wfDDs8DbZqJCtm/e5cWM76n0gG5XRb5vVSvET3qhKTbOUT3sP1tFrqSwZyT3jtqX/CvDQ0wiMWl4
HLEcYd8eu0IB4UuDbzqFQdZ4S+iu6X/jDN7jLjC38K9Jz19I1tH2WtkGSu716Zsfl3iE9a6881xZ
iRo1KXsk62PREzTS82ysR9yKrKqDsrTh4c4I/10BJoItrG7yIEaNdE4tK+0oE1WMDbkSGzCf6u5b
8plEiMBPmegePy1MUANhCEMY7X6nqDnx9tYkpVhUObTUeJ1Tn9TI4uMOuBoUOABxn2jnjjSaaHGi
UW53c3LfG+VkLPWVmjsSXvkUVmY+F7Gp3gUNk48YYdzp+v7vNIAs1JMOA79pjqLOZ6tGWTlW3zsQ
lmqyirYS9mUfV5iaV3vn765rrXEuiThbtzOxAXS8LbQo5eyjP2PgKHRW/6h2GtkSHRyadj+SudkU
NQgv2GKgi4Cy8Uo3g2gs79W2hBmZuk19QqUgoYjrY7bg/QohymACJayBzpfKs4bWRiB0jT9RJO7q
8pQc7E+6kXsHSrhE/jFPr1g2HiWo6d18Q5ECfEgiQ6nfm8kqAKCABDmhLG3mZQB6AbummPYCFxYI
Sdh2Z3mS81ZXSsWdhfKN/9XhRRqItQFEdcr78sSclNTMj7qxZaUbjooqSQUZGkZhwDQBxBuPzSC5
qZrREb/yymYE28AoPf1Tyohlg288SckKhbYXZ20QqLcJsKt+oV+ecFiW7KqY8iD2+c6RoPdlkzBr
2w6l/EnvMFF6jUUgmrBHfmwrQ3Stog6MEVrfZaydJOHQyI7FP0mLi1lT9T650dmzDOILtOaKYZ9c
lkws+0rQrkqHmOSOuy2+8FfeBeJz5h1L/L1rRd8590MihQDXcLNaarvlpsaxr7g41iDgm59FQE3K
eGPp/5kaFgjGbO/DzPWI84Z+UC/MTSujbrtO2xocH7Qz7gI82MLiumdqpDv2sqDltXRsxJjU4TcF
mYU0taXcwgFjs9kfDwQExEwhdwesRc3/cJeFPqVtzQ5OdjgyL2ejxrPufNaOaQZn2Hw0bi4j6qMU
/4S6pOVI8yJn+z5KzqHEBjJgbVfWcXRjLLvz3MMhrbP9iq0cNClmNcEFGhT7qXOVpYDSrua8WIAv
dme2d/XmS1KcNzRl1QeEMNGYDThCNTpnyviM1H+fe0gqbjffpqc3U+VuHAIW230uwraXlhEkVhqu
YrYdz41QXQT3kzxNSiZOe1Q+e881++7u1ebuyXeU9I+TCfuXi3VtdoqwPJeurwrki0mJzpZL2nSn
kkJqYPWQ2d9fMEYtBcIBIMO4toBL95jgWP0dOqOhJTrCNc1uPqk0Z62miYS64OR0UXNsi2e5ltee
wxU1DsYPYsbHklhmZr/IuSHv6g6CmV/+M3gswlQ/9dHg5eTpF4E6tTsV9YYQy52efu3C+4ImiJmu
ZcVU+kXrGF7akq0FtvodYmRSiWfUeraFbz1WxiBTmTtzy6G6O6uLp+d6K3tns4h03uDO+4R2YLlF
s3+ijs1SUC2gsiNPAmMta21JxlE5wAujXWQaAsq44qOSHUZ0iCdq8tuRNzfz7EcCkLn9bxwKyO1g
DwTsR7obAsaHih1mOzwbbzrcMsjdZ81EW4B42dWeCXriPrqjpWe2AzovXmjRDL9dfae7jicRA6Ec
ws1qdgIDvXdbADmpcbAEnRTRT8OCSxOZHdyDd4Kv0qvn7HtCbq4QBWi2LOCN9CKRJLO1bKrfPFhW
ikbPAgcF0X0d/JMOx4dTu/tRTe8Rb9PadwIL4uq+XFYSMapKB2MnljPWqtEElotHOwgjDzjClOfA
MHdAEXThZqQbUEQOBWDqxYt5K3o9QIdpPbV8t1zdzEKYZ9pZbzx2jqRUskmusjyecqjghLEkNEFL
vg1iHAqhsHxsopDd6VLxpngpJBZA1GSZRIYdq8VYBpuLXACHq21Zr8pJ0KZBvaGqFY/1pADtue3c
+I6DtLxcebOG4W3JYd3LpENtEdsm/xxEMw274uQsa1dUjAkzEwytcS12gWbHrhWa1viZQe1pW86k
dQzuI2g4sTADpAxl7Ys1dTQq6B/8UB+oQBOen1XJND0Af+OM3mRtcdcjj//6cKjZ3XpVTfuMDapf
puLvRLb6AWxBSF/pWKPvRG2lMzPv/jtJW7h4NSujJ5jxjrSTCuQHHBGBB+iH+TaukRSQCrYy4EjH
C7kkctbqyIqJ8WfWNBRR7p36k7yGG30w1iz1cOPRMCHmLgNbYyEW/AebtePt2PAMRyJZeDscGUIU
Uy6kx2t1HlxayMCP1IaLgYrtLcOc7qp8rDalP5zJd+OtJCpd29XLTUgtWcBD7ShvCBbD7yFjSiuy
LPh9mLUVs5uhy0+UcnBgcwj36FWXfPTTsV3dejJsAyQczhcOUnobuPZNeJ8lTzom03g/bjuNpZxr
SXf4uopXXCL5cMbrlAeqBdxkR4kSWCQBf3fGJX0+WVeK7i2NR7lfn1c7opsPaz0J8FmzeEka0l9O
nJg3/8dbDnPaxfqlrefhuIJE3SubFcjCEXSSQbFCrQKoAEKbDaF+7OdYI97byIVZBRlZoeFVhJa8
PJca0FGhR4j57DoYDecXEKQzJzmYTz3TZvslwYZMsACB/7cA78t2OTVOQh6ylADMZunYC8fhf+RV
gA4ILgrcS7xSenWouwS2p6nRlyvwyYSteabqTE0ETX65kYRUWDjE9UXIyTcKz+hKv7i6fKZ1DVu3
i5QaEwrwrxEgo6iiWRGx7CYPjIRpPi9I0rcwEUKAd7HGC0MLu4fb9/BDUJjW3ui0bMRlmE05iPRi
9fs7t7ByobeR6H23nD/iNyxmRNoP45D1eaZBSs4P4oJ6Cg4k1LFrZsEX9ZSVLjphVLW1C2CtfOUl
TnU5g/GYC5tbMk/dg9lPX951atvRC5o9/4TqwQ1LTBdRyiHugiJ2+0TNKlxOcyPxLjvEbGPne2MP
h8MPCxuo5sIiVl93Gu/BZLOHi+bgWi9eLhz9/0OQBqCQ3c705oU9FVxcPOMDKXIpNM5zhMOxVbbt
fqAejlvfMHk2/qgTyILMCZXWOj/zaxDpeyFBAaiKFoS05CgOZcnLk+G0Vjytgo77vzevM5rOgbNU
ZY+70TCZVupdqUvmr9MJSzPXkzp/nIqfazXs4qnjAL15iy0rg55JBF63vDr4JYiWmzsc6sVW1py1
gajU+ew5g9mw+8un9FPGwC50NkD/Gyzb/t1UNEig3Xn1mf9oOYSKUTv7n4OM3pl6E8vXWbNiiI+F
yVngl41u1UB2CH19rpps6a4FyUtCa90LhQwfyHd4pKSFxf6m4QJZ4mGASK9xq1y8l1OWwcgbj08U
Eh8m97l8+uhVkO9Gq1OUo1EYqE+hqotO7rLFqYDQz+uPY++zFop5dqXwAw4x9K6HQb99F70JBbkN
Vu0vvoklZ5jJV6TepQK27sC2WYqurq4WJn5MIY3esk8pSn+W2NHEIj9xw/s0rDW9hIuINiws5JMU
9Yt7XWc3IO3s2vVN0dusypLSGP7u3dCLxqdEy8WGIOKY95D2BqFNrne5HtwV6XS4Ntn/vYtkYzBM
eZhR3qjzUhfeenZZDUnNS83j2tmAIvmGK+x66ybgcbKaHPeK9zYGnYHkt4PFmnJFwR1GTv0fpiN4
awIrn0LwJgmm5tr1qprvCePR7e2K03FAHV5yobIlcnbRVAuEr4h9i2Sj8xqA246/R0UIJJ7SfpRt
rL7FmVtqMgynaA+tsIgSrELnZT3g0W2V+jnm1WaXs5gqVOGwr7t6laDRo6p/CrgK1s9uZmAdHHJV
0tavoV/5NtT8BKTKzVhTr+jEPXKwmQpDs0R6oY8J08lmgdfqVy1jKYFdqauvim8XsRdjxxmU36IM
RPXhZIsbMIzwVRX1sIsNBLYfY1HG5PVBBSTKolxJ78zSnH8SaWpJbJRbbvurqrIgbHeo/Ypq4XKU
81E1A39Dy+SVSrpOSQIXPbbeveWuZ4wYbWR3+v5dIK7znmR52d/sbXFOA1q0Ov/tkXfjwKyL0uYH
jAYQWAIgR99pBgYTl8ypUTBOR6xVzgmByqHXUBxZ8kjoiRS81EPvJ13QX/DTytkYfUWs0VFFeLta
n/R0Iqbk25PqQdsNqSPkuPxR++4C3uhP/QDnoWyeyTX7L8eiMGnImvCdy4SxPq9+NI5v+y8HoVqT
FTMv+vNbb3Fyh8W2/G5514Kw8gV7D7aWXT/E4iaf1t3ScffPh+CihFWE2yQwx2XS2WkvI4Yj+7bq
38Seje3S6gWqezMjt40muxv9uFiXlVfydMCRk2/hX0P0j+Ss83SWBkqmhdvP88fPuwTNKT3VPZip
vSwCuvPqPWfb9g/W3R32kWh/ZEzFXzMzTGkPOjhHg43Y9dM4++g81P08YqJiJVkxVCy7m6H9AijX
Im0ak/eOAvgfmtoKs5jO2hNOgcfIpM9irSbYNMIn9Uo+QYVgXBxfZxkEoRvRaYVvp4H+qim6xdzz
a/YKMizzkpCyPKzNbjorsCCXfqDlYyul2jvs5/7Lrzo/8K649cHSXamF4rC0VQ8HsdyCnFyykhpR
sCGrq3SmhayXU/836eN6IvGaRneNDxugbA8a4MtEdXQsFBTWzCJl7PiBad5PqxhEO1zHrF+WKWqi
9kPTP54g3aN/a0eBZDDvGogPYURjiL9ZfIlQahv6X2iYLUNilQ5g9xEfqdB9W+yjKjggCi7buiSF
E64dAWGw/0zmqB2Ee7l7eexXGFP7CQ35Zf/RbzLL7hRN+szAvZ9UOq2OFtHy6hpXcZ4G4GHwvw0R
zO3OG6oDBStEBxX/7dwj1Ziwk2pzci7bw9Ix0OuRq7AgUXSdEz7B8LkaoIbQ+L1sK6BFHivwKSH2
Z946Z1IdjbXJaRBAqNGEZOzzPeF1j0E1y6tQKwKZHagSAYe6rCsqe9wbn1/TKoF8IjA3K4cb/d/G
TLTvG8R9sjSBz8qwTzzpLsaAcLnGdSbZFsa/BqIyFKRrJuQbQwrR/hoEKKvmzLMm+wiMNV7lWrCY
tpRVNXPGAxj6wfAtGM9cdNSAyFjY+3aGaA36zxIwRymwgEKUrDaymtP0AaW9VRyQPtkaseAdUaDg
xtaPrPWOawoOWGctoyjb/ZdpUS7pbh84I6YgLl9rr18xyP7Vd8J+kosg0b/rJm5WnXYcAuLfMBik
OYrwYxI6B6nxRhJkNWdmb7RilnmKEhWi+dOcj5fKAzemeh/whA+i7uVT380oc13Tc7Teg09aLAWT
ORxojOAhQl1ttZkaxXdgAOUsFzDw8xCuaDm/c/6dwYfOKAad7LJ/XT9QZs3pBhcxpVRSQNGUSoNw
Ahfdj406THlcYaD5RQrAjjZbSj4zTwYzL7K0t20oBWSizCrfD4UV9m1cgEmleKwyRgi2QM4BL7UZ
N+S6gtuhDxwPMLQ3GpAZeYvB7n0Hdgsmk/0Bf5F/09Ywjkqd104seVQii5PAFzbCdXRY6NrljIuO
a1U5aed85IE2RQ+nXNu/d00SKelSxklZOy1+qYjwRJLYIUVD3ATY/PTiKqfv0ukIkRpDwQICBZK1
YxV3cVtkWb4ZRTrFT/mYcTO8ZESYMab1B23eOxRHnO+wYUEtmQcTkh+zbyAapQANiSirsnZ2PD5q
gJhP0ClejbzybvAJsVJF10NpXpHK/KzkJXsN6i/EqdI9bS0p/cXnjyv2y2ONNY9Ru2Fnjr/TaZUw
bx2FychvpTTy/2EiKsL0GwXysTZ1WdI4uDEeX8+ELGJX55+v2IPeS+sNCl+aLiNe6BbLRGChHsqK
c0udaIO4s/nx4jUu6RXJcKXOzsPPzFxyM3+YXKt9/KCNN+Adzh7Lqb9HdRcgff8KrqbHTnJAXoC3
nVae2ULaDWEK64yWXimo1r+t2aKLtlkB2V2nM1YS1dG+lyWYTQE6WPUvbrOsuFCWlNrB+xPaXZt+
78RIrT7r/aBcFJE/4ijXcM22Ey0qgN+IqsnJRjfnd1+BBLlE90/CSXJK7wn7OTYIkY53Ick7Q5d+
VDNm1X38nD+pVTG8eQ7urDDq2xfg/lTHNKMCnSkHLg5KT2leDJkiqDTxtAsv6okeO8A+1WWpjvDq
N0mfctIdqaIsbaobfixBmeQQ0dETHVD/gLkg5c9n5Z/fmhd1N+a5kha7FNNz28DaXk2rHvthVp3R
vW4ese00s5jtVadqLNfBgWjm9vyzK4jS+dFnq1A5oYW5TjAg/eFa+nXWbFf46WJM6gX569aDDxX8
uZfWPMhopXyac5teo9KvVMDyliVpJyQ+F9zGEKCNCDcXjVnW5rpCZQqYQmiSC+IwY6BmYHs1zIxg
1XPAfIvn4QrFxqsd2Q4TZc7CK4d9PbjuC6POLYJRaN8Li3jQD58S32wvVogPTqBZ98FVIpasW+9r
VlCUm/HvbKoC1FAcWvojJjpiHF0I5eBDnuDgT0neOK9NLyyslAIQNXdSdvgClCJtRHvE4oqgD4bC
N75dfzJ5RqO/FFzl3mNDfaw/+/R/KuXcrfWvUMwHQeQBqFzfsM57pAmdlfImzImV2/iZr7NR0XVd
IqB54kYX9pJ/hi+cnpnmm2zqvGQMsw3u9JGAI6WxhalmHVnwsOdDim6Tia8koQaf95FDeLH6fhgw
pl6KoOV9tjkbyMIZ0qaR4o2GOrfaMe3iRYfvdNzj73uAHZEpUbdeeZMzQ2hS9Kv0zUCD6xAF3nHU
3zL1INRkSxFVX7ZTigRUdz19nCvClw4+t2ZDDegLs9zefYzmu+1gDFw1HlcbDwidG4jL/zWnqJFr
hKcsAUoUUOq8Rf1sFBol9ilL6qhIUewgabZJ/E0IT9cwVPOMwfIgF9dT38fuisKlACnYiR5pczs8
XB/xeT04Csh5h0RZRZ/+AHzCxZ7mZ442vz/sTWU+thPp+kkaxGWNeXwyki5xx3OODBVFaymLNQ69
HfwHmc7fv9OtSIcfOSBAbdEK1RRSWx/Ao9vn6hkcrN183teqTX1ru8kv0alS08vUIQ0+vHfzkTws
GMH88+NanuvLhQkJt3cHFtNnjr9Gzb0aYgQaJ07xcF2rhJOxLlfaxvBJyTf5EN8/GdifCXgA2gpY
qeU/GaAfMHAxpKPIl0NROM0hPdBSCoxjLE1pjun8yWE2NWHJ0CmS4kq5iP2qhTj7xJSt9XFQIvNA
OL/DZham3P01xvWqdTJS9aPHkEVaFyMbx/vN2y5vwiJ3AJH8f6tGq9hoBicwSqXtlxRqN9T+pkZ/
E8FUNBK4/NSTz6qwq+WZ2U5mXfeyfmoeZSG2hxypw63PlqETSX+CTbbqAOhGgVHOxOlU0NVN5E9x
jf6P3RmulLN3tWVa4XP4wiwy7o0FHy0w9g7MzEigVk3B/3vVHZe+7VRDNYzYbIfpmZEJipSYGESQ
50J/NXAmRsRFCOg81VznjxUg3nMLvnk51j7lpLGJ/GkCdHkFz3uWxqFL8ERTgHibU8ANfyInv0hM
f+ntQUm7+b4lPuu0F4R95jzuTbt9oWTVDYzUbcbEhQo2qn2lOY79ysFWsSEp8hPb5pC2YuOK250f
8sUwIlmqEoqkLygDVlbJZvc/pFPSYOt37MtukeXdrsNZGhTLkUVAz9v2h6Td0CzDJZ0SDjHWxanY
82YDXoY2RQAG3dmbP2w7HLV4FR1AZ0PWGElYNRIL/XmSe3uU4IfZ6faygnsLpUVc5Vb4/M/SJt4D
+Nnszq/eTUcVMFppbSy1uLM5B2wFADG3QFXiCWV2kJkTovgkYiKkxtyH2HKBgNJtv4lRR9k/aWCS
pJwiOML4ehcqsLr4G+oadF7JCj3RqB1BO7vQJn9ZyE67NOyddKgtiUr20ksv7huxNwHI5xlu9RJk
5LRprsTIuAEZXHkg0n+8wRTeWSI2ecXlxnaUflI0Xu4k87OA/JJlDlMv7/kDUUlydijvIqwtVY+S
U+mOgTpEpRPdzRoeYN8shYWtl36rJE8LeExBisvN/OJtO9r3Qw5Ml3jAANkSsYJS2lSdc68fRtr8
KT1PWgkzzUpfezTwcfioMAYKzXaUyv5kPa2K5ieGXlqrdFWW4ZeHBXl3TY0FjZDTW0iEjY4v4S00
6djp7RjCmanSrfo6Uk+sqIBRKjlYHiEn7ky2oaZBqabOZDV7CtPHCP5oMNgh5oL1JHWy2T5QrtPz
B3w5VchycjQ0QFoRSLAq4fn4I+nqIE0DOtXOJzepaI8tNKGIaxYQi+L+Oy5G8U4VW2kMmVT+cV8N
nRbaBl3e6+a3QRaPeTfun3i1S5skZdzyrZMGMSA81fdrunfd7xDdhNzTIcCbq0ILH5+t5gB5auvO
S1nH0THdfXzCyXn3EBzKq0nFy7layFiD14lhDtv3IlnTIQuXhoQHXQRKCyALWknB5KYdfaBsEzIJ
3P/7SvozcdwWP2xNCITlpG2YjOitp6Z+4QkThcAhcGXincoXVP9vMtg9dGplwGZ9uhjRnCzBWJVG
gS8hcbvP/sQtX5QIbFITbvytRNZH9Fk1X9apoTmvYE71gd3p6XtyaqdDQzSCdgujhDaVQrTBzG5d
MKcRYRQ09rhkB/vO0HxElK2qCDV6GGEmM09uDltTfSvDs2Mo4lYFkoAeqYLRrKrZOiJFGaGqebVk
ERt8uDBz7HtLoocUkVMfvmwBkdkkg92ENX0EOFRyChufr9c4FTTB/CNX/4rpR0xUpNAMoVY0z7qo
TiJYe4mM1LAFiuW+hDvsYiM+PcgZzoCcX1Y5cx/6AWJgssNVuiCCHljbWkjIHzW4gUtqKNkfxEiI
h+JpVeyioEdGHRU8UsxTbBD1MNhu5IGziGXtB+8GhHRWsNQiR145SO/tUMXCAcg/i0qiN+faF7Ir
R2VVEoRJARRo8HbnyuauSnZdL6mZLWYOBWE2CQr33qLZ5t2bMe/Hx+uloHKpzzDNARkvKrCIqCkF
/7F4Qh7l51uq/81TJDuBgWqMKzQ1LLBHCW8RaURG1qwy4fXh47JGza8zAhHwMNorpjrlgCL0W9s+
DA5jifd8/1NTjNeQgkyBzNk8h/YIn5c2/ph0TSCgziK8SnSX7fOm60/p2v5lFYmMkl8ugaeMsC2P
jmn1Q+TTkVkHd+IhGDglKPllbyas/3nqj8clHR/C/pkQyHZkzzN06QPu+0TOOBY5dgAi1EQ2dVjL
gxE/lP7fj0VYtdwyLq9vOfViDECcvWuXb1NrHkOyMNA33Ii5kUcqgqcl8/HGdDdeyh6hYHVgQ1iU
5DMhH/kFq/WfdKVqpJybVxfAlzBQEwohxpS5yP3b6MPPVIaZTiTMKcOR2ABZ2vM1u4lvkck9/gxL
ayNZrRZnCD3I9us0gIxLpdAOmt4s96wPfREhApec1dWJ0RRtiIYo1iY2zN9m1azFhAPJfdKK28ZU
cooqWDX+PdjiYbDwnQIj6F+RHg3ssRoOaOkRllC7Gk8bvxHUCA+zQXHCaE+tU9WzinVRWwd1U7ty
Hd2bZ/jrFvYfEgiT4Lbouw2ncUIaYp6bbfNCnvmLcF0BX6BE5UMwohMKrUhIxz818rNoRGd3ZJSy
sDF+ZdVBWNgNfW/jBYRU/RL4zlZFzdMNqI38aQTlLoh4TTjDq1o4z2Na++nh2Fg7m7ZLbdGKwwgy
iNm8WU87amn+jK9yaUI9ZoAWCD/6mtySHfddb/TTnYKG6/W2/FDMjrMH9/7EJI9jcz4sFwAKRZaJ
IF6pVKqu2mEvlahw+n87BnTOLd6VGpCBC4FybfnevfBBOB1MVeUGYMRXqY2fiwv+K7t01jsR7izb
J8+/DuQhWzeZiZS+B+I4WjmGyffhYQsbtb8G5gzWDj3Fx3SQScFmdIIOshccGBBqEN0EpSTqRMJa
/BeSNDnQC6EK8+BJHDegq5E2CpbMFs3AB42rg8L059O8y7R8qIMywB+jv/Ae/QIuFuQvFQ/1IXLd
xSpJpSuzLxUh7/dnM+KvQgWO4nezAFXAA1Wu2W6CKxy6O71Mg7XOZO6kwizMUWbuoz9/CxLujDgP
NcGMQigM8N6fiQg6wZEDea2RG6vKH4xidKyy/VMq5G0duphyr8LDiK9pEa7is1a8U40lrhdrrL1G
1tB1Ww8leAAN5mph4+Si2Rh6K1JQPIzf7TGfnm9Bbc5Ocukbi56nDmR7bO3TrnNUobjWIndwq//z
CZSvgOWc/BmpA4k3DsCzAyygJ2nHGxxxfiQ0uMRMutWkxJ/sulJgQBCp7MW5gjoYM7RF5z7GTZ97
kS+PgNl+ruYTj33xqNiX4l1TwkpbP2dB+fdwCUO/vEEmveQvSByWP1jmyBRipXy91eaSLdgF+fEg
vK5UGzZH7jc/CN1b3f8hUVPNe/Sq0zo8uC3m/jc4Ywdn+JOgd0FHLxJz00z6gDE4hdR0YBFVZ3ED
IDej05lJ3phRMr0HrpgxE4Uets+jz+o3mS4ESC6UHd2Am0p7nMlovrQDpulJTyTUhTCkdlJ9+oKt
5V8oL9virnvFI4qtUTwZgXYqllr/REWeLgizNvPe8vGnNlr6p4nKVMSA3FpgpoNuNK51GcER17WN
+w+LTvQsBggFY8swqz1NQwDPP3Jk2a/35Y4vdZRl9NYD8VT7+eJ+nRQS6dw3L0BSphRwf1j7TXOp
rBcARSViZ8mtOiegOTC47bMA2K35C1MA6jb8QEpVpgaPvpC2nLjYFJbiGz5msqFNJAwn/2k/FOTw
2U+XjFHS6Uht2giRINC8Y8lip27+GjW736ijTdCPzCIo4ttnOf2M0tHd+JIhECfTB5pOCYk6tPIZ
4Pk1Tu4J0DMtexb9oj+TtAYd6cXSKl0lfEbBuEgtV/gRbXbFZWtpckhATb2fTmF62HAfA2nnbE1x
+gdtdyG3cmGj/uxPCubrz7fIBP/gwlOb1Cjfap1aYN/VqNAtZ9imMh56ji/m4JYvAHiFE8/uLXtS
I6BddPABRLti2GDTxWtOOPXCs3JR9II5tYuMJs3/+LXnQ4wOhtJtsuTLqKqSyIC/f03gofoSza2R
zLdb3t+SCXboM1pkZ8SHf72CkC0xFHWkIPRDLlIGJEZjEv6aLc7MCDO/BHWVck33EN7UncCo4W0a
Bsd9VlpJhJZWC9NIpFSEZFrpd33+fzt81FOZVyjxk5OR2y1exdDqlOKxBokuTKZcGhqefVUbSr7J
YE818iro/t/1OkqVnsJuIjBu2MPY5FnFEkopX85Z22AMMauXWTaDR//m3zs5HHP65ffUlLQAKyWj
ClrwcT9wNKUKRxWCQeSMByHHXTi4ttVmuZGkvBMUpqDh38MiMunBbnaGd+mnSkE3NmjLFLQy+qqz
y7aQo+ysSRjHxngLS64ZASC0xY63GSjg0d1zRVV1NjPVW1h09/o0fmI7onLvbrVo58lBHuP5E/eF
81QpfR0NVI7Bu6Vnq7AfN8gIY+kQOA6zz+PQfsIsmF1QbrrV5WeKqv9wT6ybwBlMcvG+4mtvI549
DcVOZnlpYpZC/nPk/JiSxyrroZFHD3TVMhCxrTfv3cVmEE9UD4V5GsKI4BI3feCBRDklD6i/VUDW
4yI6zes/mVzEPog6aKj3FOBujuERV04gpTo4FpLLEWWWix9K2ABrMpzV8sPtDlUdR0XNBtTlFtvn
iiAbto+eOR7wnzo1Rj4lid1p5xpGB+CHIgtFgsLIhvHPKfdXXMW5JqiDTQbpkN4APCFXYesX8pwz
1JMKFvjq5ONj7IH5Z2pUrfx+d6rURffl9/FRjXvHfSpVF3vVchLmJasObbvAkppTt2h7w77BISLl
WpoB8clWKijgD2foyL9OBJ8rNLRKslhxdiZwLq+B5vjGnV35IVXKFNUAdUzKoasEO0kqzBfBrJq/
JwcZ90AUrb9xvfDRvLTutLBHf0w/ejET4nUGUriYszL6nQDEKQX/FtaLCA5wG3N+4t1oBC0ZCsr/
Rhd9dibQFXuDPC8evJNp+YwM9CWdbp0/Lf/s/BdLGhoyxIN+7qHH+BJ/jBz5Im3I8RlQgktMoydL
HIX06pwOeKtidviCcVVyMFl6RD0X7/hHp7Su/sCJ3mdv0E9OsQpbbxVroXAiZmxrclDDA3qdYOcm
xsbl5v0jI+tGSSaqmuoEkl5T2rOFekkMT4fyvq60WnEm6VY4E6lfHOpmnBm/qX23+T49V/4z6eaG
5Q97ob9euAXkHAla1e0q2GYCYHPvAHft2fpa+aSbEIPTKPrVAfWY6GjJGCGEVCjTtz4ld7g5/WhR
fOO7ZzT24OpPoxvYjBm0pfUd2YTXH5ff0T9XmLAVQ32CCyn+FlLEhZrStrPCENj+Lxexbl1zfh9I
YqWpXiny3PBDy3FjG9gPzibMZFbtKNwBQyBAmfjPXpctFpd4hTanRcyIwvHlTd316ufDjb4lMJTc
dFLY06wrU0YU0JI0hEvJd6REuFXyNLOsrsbx3Uekp1xj71fxjmCpnQaZCWgjN+iNcMpVBs7jOTIx
UfxD20eNzbPDNyvbmPD2kRhw0FlfN6/0+brDS3hzD20jLyFqnOPbOexVubLRVCACcDM3yanlym3/
xEOi6m3K5vlG+f+gW48EHmEXl/sZHl7vPm/bmgbNWsfwFb1DUVo7vNLR41/9za1HQhFl1IIAaVPM
sWiV4/EwLjEyxE2GWvhjXiyt8r8iqBMgUkeWDyYL9m9j8PijcvQdbuMN6T6aNfdGHb8gh4NYfX03
VWRadJEqqgOyAQ6C89GVCJGwZ/ttnkCqgUU0B5cl3JQEMUiOz0DUdma2N92bYngm+DEPU47z83AG
Ssx/5AhEedruUojWnFsOLkUXzcExuz6EwmRmngfJ8DZmUqDV9NI5DpE+s9hgSU8MAFc8tMimJ7yp
LyFACNhgNvbi+3+4tVDAc1RYHQd8VeeYR900I9lUM3Es4+obWUtd42IDL69o9zubEwJUTLwRKPJe
vrftPhHb0VYsiUfyICRwT6jKpqbZNNNQAG5NVoQoLRjkRLPXK9NuAG/D8k6r6OnQFhmZkDvQ9B6h
A8DgshUcX0HHTGr16cxPyg0JdTCqUCyeTjwaHevaByPbDC7xZevj9RSE/UgHO1ZeEzfb/CPEN1Dl
+sG4EN6iOWfGauofULKnt2r1Sqw+3j2oaNJ+eQY9ubNxR63U19x0tsokRzaFeJrFBFTkzOtGQOJm
dgvNwcjxMwEzSEieAvd1vaUfQ+w2vRt71V6GXa9KU3iP2iSYlr+XP/wVJiDHtux+MVk3RO76KWez
UMzDibcJBdRGz1URPtXyuhTiPa0aJ638QEPpHD1L1PHt3vdQt5aHNcYWj+fOEV293tqfBXMEhdU0
7PRl/1fpM2kGsM1rRKIpmHB8VOOVmtQK6O3OO21k89r+1ebnFyj3/cQ/JlkWGHyfmUkYfYwMdyGt
W4zS4ZByL+XYl0pQKEO4lvcEbqz/rAutMSMr6cdwVQUmyQBXSJB9rHWuh9yG1P5e/oS38TvwAYYO
iYTAextXnISuQBL+wBzrWl42nxKBA54sH9x4OPWobdNr+rcduDhyGNU+6xXB2imLhuetbGjv/prM
/NyAIm3NZleJBYgKEloFTTmEq5AX8VuhVFoPQ9t+8GPjT8JCEGlLlp8qSXNJIVyVdlxKkD3pQ8YQ
MlQJn1s4IIEaFxcRHN+HDbXswC0WCUdkfxeERiWNPY9XkyatpwYl264nM1gVDc+bklXEIZAUN+YC
IB9ZGulsJVDj818TlQD1aQ6wxqxgAfc0s7rZ33i8zStxadNPoY5lUEBghm4ST/MHLnA2k0WxMNse
jbl+9/3Hct9kFWiubHhRe+J1yBLwN4m59AtlwF6LuSGhYUsoqDewQ83CzT1IPITGWdy/VlnwcCGE
pmGxwQ9oBpDRkHsEEb8ONg36KM08htWd0vmCbrk+GNK2wmCYrVdhGjkijbZhGHsP83h4IHkFoXpg
y+9svWsqKC350tp1E6UZfm3bIkbWgPhSjSxqPaOiIWCpVY+veZhNCUFaYE2CC7NOloIaiS9sgDzA
o/Tg7jWlVwLeHjkEOg2yEcYKuTcSlyepz/6ZgCcPgAjCDlCZvYsO1Z862SjIsMZVIr0wiaTTd05p
2RncIQ/VbtY2LC/Uwjq/5BJSWQdzLDU7JP8kVbAcWqCGk2f6D5k8nibyA7yGTTetJ4vaJ5YTwv9K
jhq95fGxDimHMje1Ou1uaK6ZBJCnlCE5aQP6iZBxuUQF4IY0lan//IfD7pnygR9dcMXWp4NCvtFa
UwEK6oVetvSPoqsKaxSrUzgwVfTyLMQ0OFwFaSyB1uAIfcnf9Tzsc1QjNWioA+cMZT5xaXh/k9q2
+lFAwGtjle3/7FATAQHf44k8EJyH2t4QuqGjtNiQW7LmA2rVc15OBPobVdMYEWixYt8lMYbgXgWe
88JBwkPB6Z07vf+bXP/9VntKu8qIBernu6xOEGA1MKDtrIky9aMRVImqHmFdVqCqi4iK8sVl8Wo7
04jF6QiZNFMYpvgymE7UBR/jv2UfIhE4VM7DdjO6mnvdmGhYqnbsHbbpyWXKgw4SuWhsE1V1Kd8q
sScOBkiqSGoWGoBvhMQneNU2Cy70qZ2e5cGG+TbSdbgaRrWQxpSs9SwnUWwYDJ30jdDBpzZTtgZ/
Iygs59NxrarWo2nPaB/xVC5y45G0frH8wpruQfoibUAdsh3j937xjBABhkfMPY7erch0Gon49tw/
hu/Xb3I9NCwr7JJkkxe9J1Z9lVyIUjA9GRGxo4/nZV0sv2BPL2NYfpXy82OkmvQnvxNUBLqkvgwW
KzfBIahYraOwXJRNePZU7la1ouBHBBp2OHND4dQfTjYg/W9T7HMD2EWGWhhOohMHGzRJ5oBhVTuf
uhazvlUalVuLSadAbLtJYCApjE1ZLzO8XvyeOpRtNr1EinUBTUP/3UITY3jOHjYM87ibCCNubxwa
Wa31xVnSfXulw/GigvBUf4cznTKRCfeCad/RehMpKEHalwGchqx7ZzDV8xDza/3X1Q/9nLfN6u+K
jckrDPwzxGLifSd5619EKDQz31xUuU1FS4aOAoauKnmJSq/yxbJM7ahy8rJztVO9O6j1t09DkOg2
X7H8BcrTb7dbXh9W5GLmf6+d9E2nxVqVG/eJCiFwPCAsHoE3rr3/BfBwaxWDlsvpf5yAT01INg92
Zo196fF8SabjzK3ZV30ua97/Pucd8wx/pVpurldR0EUI4kyg1a3nt0o4qu3tf7FF0+AXHIEoHlqE
jd+qjTVEHP9s1frZZEsLiB06NApZ9hv0A9HWAdEopUj74P5EfGs2F3QPGG/krIFhix+JyjenNq47
ELL1K2GsdVlJj0UncDhbD/qgMUiEX+bHkZjHi/5kYRTQqbl56AxBh3jPZHCzD77Hu9bJD4VqotrJ
Obcl5TZe9TDSJcoxCFzJfewdY/hGa/+7UhZeR8xEZpFUGMVyzX544wwXxGhtX55bkGYvN0ud2Xx+
+N8lQxImXinmPDDCeUV0w45p+s0g93Igu1QiZsZGXHi/Xie9PO4CPf2pyV3UEPTOkVEm1RB4ZmWT
iIlcruq9lh4DrO0U9GwOyM+vOej6QkFtXcVMSvPAC6H9XcHRrhM//cWhMKLxezbD6UDZz9gEptP0
Q3VaYnINasAJk6NbWus4d8GNjf93Rd/FP8nZ/q5fFWajnC8Zmj0j+PnP6oRlEpC06gfqgH7GeeM6
AHQCSzDLGbvFKlnJHjUGhmLDO9LPFvJjqZ5QHiY+geN0fiabqUFORJlYWjuwpLzRg/EL/8VsCLEn
H7CD1VBdclbXvEPjzHgS4cfeZ1EeMnJdUsUHy2VhAMWE0nzX+F4/CYgO8KZRSvav4oqLy4soeabF
IVmLeOcNMRKNLe+wJm1Mw4Nw0zBd4PLwfCsglzfXOOvTDKSIQIT3DIqiXeyjV8IxcXEDYlXsiTOZ
12PTqrRGo96KEGzAdqgNg6N+daYNLklOYAop7YFbeiY1l/zk/WBKvWZVBNWE4CRcIGXPjfcbQ2FQ
AZ5Om38XmO7LSq7lg14HSPGHkAjCUVTUQ5KLZI/kA48AWKo+exxva8feDHh48AiQVRLRoZS3prFL
VqbWRcj3m3eh+5j/ECjIvFC6Q0oWNIEB1AWALO0vLzB6JZq8TnLNEYJ5avtjf7SKtNZiIq2qv3vS
DDvkthN2vUtgOWhVC1fEROLHKw1EgQTwyzUmC9b1jl0rjWtoupf3Q5yGZ2UqlSHmucJ/uAGft//x
KmkuiNXu3r3qm5cg/3YZMiUvPK7pXPdjFBGe+yR/qVe0kSfRo2kPT/Om8J28RZtr96HDRZFv2vK+
nBi4CWmmXsBzsjIMMsCU3qVhtegIhPKVrBLZ25JATzLiJXYt+RvUnYFuULJQYRrLWPO/YBW2G9rX
iY0OlaVxXu4FwuMw/1zviqUf1T4LPrc2x09WkMT3qfD53Lt2iNVtHkt7F8DgP4G3ojLVEYaOrLcC
NtYLn7kVtdMwhi3Uwlck04Pm9Qq5xuMWKYCg2xRBTBmJT10eY3mpw5pUFndNqiZo2WQDYKAjoK92
OFv4LOPdczgW5gfTaGd85x5EqFHBuMXWPBJvqdaf6YJIX93MHO5o/QQrXFW2OVscitKU+ft/1mYN
W0rl/iif4uR5BKbbGKNRcDOPB0mx6QKGB1AkuXmypb5Sg6KwXrMIAXkaHujJrEB0AHpucuug3KsL
xiTIJNl9u5MG7+yPhiPc4EOGLKSdhujK8oxW0LLR2pKZyA/9HV5Hgccwzg5H5iG23YYM+4Mp9dZE
Sp2/nhxgpLL90uY1eChuO9nr03Es+d0u79hyBuYfsIDuhjIOf4UJu6+lFR0s210KnJH3Ig7CAXSD
b7DIhm01vMZ1Ug1g2VXWGPodcWqTdk1Dk25yWjsH3+I0Au2hXQlFO2m0kJ78u5dw67qGdUdOeOuJ
0BpcCecHLv6KS+viQ4iQeCzEpzKDvgPduhZU0q8sh94nHYVBs929sp/UcyJIUzL5IH+c4HW7nenP
+yBCxLCLJuJ4RynE+B48tOYl1DBaZ1L1btwq72PgJ8UovU/rXr6pC9a7uKEsWcDu41+mZrU/vp8h
BCoR/bou7wim8ic7eH0HHhx6twZV8LuW1bpv1+RFmrJHZOwopNcaEHhpoVwi345RmGKnuLBw6rAd
IOVcgxhEQXwFiCWbGApz+MBA9tkab7/N3/9Lliq8WpCFMLQr1M4wC4vyiO/niFTDuIOuIU6gHqks
LkiQNa7ZpYSj9OFJo3kFsQ2otTeq/kEydAobG62Q/90DsmKRxJ8zx9EKvfd2lUqxbCnFFgTi/mVn
s/jiSTEOgxmeW8gQ+u1oIBg2IGhf3Dy9neXPRKbha4sI4ZbK0zdk6PKNMlRCu03kXtT2bG1i6VrH
VbxRgANsaWvnlK8ScVIYG6NffAvK/FVgl+qNn/fxR2AZH3fX0MbLM42Lbyx74Z5EyW2UyHxLLyzl
3JwBLXTNy3ifsvO0i67tk3iCRvqyGQIjff2t/JqCjegV+WsiiMTivmo93jV48+hVQU5fSompbCt+
MDkdQBC+MZPcJaJaOi4epeKybEVktcFVpSO128wiOT5ykSNeBshrS8KuBjjopmLOHyznH1v0KI7/
FDoazF5djBg2fV00Az/uBFxbyy1m4vx+bRc0JsQgMLkfgkaoaKKREDW8ACt0J/0nWOckDWA7Y7JQ
mSROJrzqXqVWF/F3Wa8GtXK+5TMG5rHISRYTQaSmu9Yem/ds7N0biivwSTZVUSANHFlPc192KWcE
23CmxNe6SQ6f5tYPRZPfyU/PBXgaiO2rmotKQ8nvkqefGSxsFbkYTJBuTSAfVwf0gpTYMRqoE8tH
zP8OsrYBvRD4GwO/ma2+JDeTUt3dAXtihAzVkDXBYOkwn7gfLZNn8p1T3MkIXXAb1lwMbHi5lPlh
BsnIGb/WmD3pQNkuNuCkbRi9c77WynT1Ylhbr0RDZDgsIA7ID+zW7AhBndF9DiqILWm2ym/1rJFD
vc3LqKNNCH99imHkh5eeE4G7MTC+y2+bTRXtKYk8e+cqSOxQT+dNs1BOOa5fbX9zsrRqBV9lgZwH
yKVq8QmdUNEuhNhAcgoWwPXs7jvJwSlbleCgxsFiPIO25CgxYS70lOTgff1w4MLkqgYkOmJVkU4d
+tZ2XxXGUw+D24SD8KLR6iXMriw45LLV5KoP1bT/XEi2uxLvWDYZYmjCPwJqBY5I56TxOiYKOKb1
sItGGgaau6JV0qOo50KOfxHUB7HGDmAZpx1J/stSh1PoCMDUbtAr0OPSzgdfIgf4fgKwqexbCe+h
OZOMaQNSwlKuw44CnjbTmqylsHn/v4p3JyWst2W+Lp/cMNyVPidA817Szzh1dYKf6slk7PMBMaH9
MMOQBukE/TaQhIfyftiGUJikaKXyYsotRyg6tKJkgura90RVJBM4TqKf1HAqg3K5uWktMeSaQ9e4
BBIC7Xodo0+lSKFtDPbDoE/OV59GocngKBGjRg6vaCzCVxCOhWuy1BlAoYR8R7zmbivkgvmkloyZ
FC8wEznhFUKGXZLcYWhZAbxOa+3KgWqPD/TD1Kv8JLxtbqoJZ65MsY+NTDRbEGI2/fMX205UkXiG
MkUrok5clo4mz9EW9ImE7lPhjeRlAFzTVn83YrWPjnU655B/vUY7opdJrR7tO2Zwlxfnm+wYcJkV
8CCLIUu0GL4E8qHjYJLDBk/RPG2/bnEJgXIyn8E/RGAgCIobmyyR1zuvr9y7jTFNxXh1ozFhEN2r
NYdXkkT4XzTMrl6Tg9BHev8DoClU7aiTnmPPhkLmBjjuu3XFZpclnVnmOxGUWAGqZafF4t63cndq
poiKIyi2Uh8/0Dvg1VauF+S/SnAmymdUYk4/z8/mizoXEb4CjkULayLDfKYOo8NRpkJ4B1XOrT9B
dqtbChBvt92AhuYKMfTRFvb/e4yrLT+pLdio+dzID4xHHjsc6oO5/G+B9peEg4dYNGJr58xvEEVs
hnWI4SJ6783WNCRYCU3C6Vcojr5mn4Nk0zt7VAxolW5AjKwRLaVFHrprcHONAk8HTjeSLp/bRnp4
smXJIwzp4vhx4CNfCaI9W3zYLK2cFhCWLyJdeLIhxqrLYUHz1vG8WkRsZJn17dyttWdaFAAmB1+p
USMEgjGlFfaV5OtQsT56SVCnTY6JRoZhSAixOi7OxdT3U6iTph8aEIScTrm5QQcpijA1E3wHxJ8k
3IRss3dSzLBQ+5CO7yDccAaY+GE528GKnKk1Fv4S84i5jhoF49cKm4ozav6DBtdC1ivvbMn2pnFi
hKtItCKvGdhg7kHMiuU7Lsc681xPtH7lVuS86xPKE3h9ziX6m2iQ4UtFhZCbetpaG6sYJ+H0o8Vp
O2ocx6BqS/GkW0Z1KqPze7wYxhxvghW69avSIL7s1EiDutm8t/U3MhacWwUQj9jYI0JfujxM8g4a
iSqM2Tc5eCRqEW91U9yXpP+LAOQHXBpAFo413kIZ6btWHgX8iWk5gmrSTVA/JUV+X2E/s4Ks+REJ
2FJQMp7DlPjK5MYUVfYEUiIcLYiVtQVEAS4cR9nnjFllszCU/d6fzldD2V0lbz3afNByNvyYWKOn
/PvHG1upE6b00kU4uoxSTaZ72zCr7FAeh8Ml4PK6g6zKwNpjM9uc+KT1n1T8n0ASqUJX+iOqQvSR
oKPMYfFkWpuD6jhdmYQ4oOcvxxX7lT84JJHlB6Fl9Y9U9Q/cpdzDH9vYge3RfTZ6Xc8Hz5cWqH2R
RJWYsXH926kYXB1ndFz/lWzc5jGgjOE4npRN+bsT5KT03+zkHPgU+rPPGJ6ozQFX52F23FZmjt/T
jDAF5iTYtfk+wc/HwJ42gb1n0aZpJ400rt/c6f9Rdrd9G9o43gFwmtAlpwvyFSASMlBvliNh3pcW
MbYOvIczsWqgkdg6fco59HNrxbhh5hyGROysLhFGBCKIwJ+fn3mVofr0UI00Xx7/+KV4arQlh8WY
VlRQsi7IRcGEBfQYiZcrNsMtV+E/fPN4QR7p19dSwC6w4IVWLn8dpg8Pibj3YeMDob4nNPW3Sl8Q
wkpCEWQw4Lc5PV74NX0Wk1+mL2ep6suEoHXWon4Y8H6XGpZ7ok3IH7WO9lXSLMJyzLQAz7g13BL9
vnu7Yr9in19z/Hu03DLbVI5UJGCROm4zeDrNagO/7Kjwaet//7fgZ8g25SJdvolgX2SxzzM3YFvh
Bm7HzGsNRWULoJH2dqnkb05jtlLZGudpWPk1HBlpH7eSnq7lhZK62srp3Z3gSx093YdjNx/43Cpp
bUiQjVa19QN6xk/JwaA50tXYy00zrZyEkW1jQfRtcGhr7rsVIpO6Z8Rks5kA1EvMvjmUmYB1ABdZ
2tReTJ0evrAGSH1qoiMPzK0gLq9/zyJNjQcI+bj1remhxMVMkzzLg6x0HSyt0e8dj1ONt15efBxU
Rw7ZIxTcRhv7K7gVdTOQA9s5Jn24+RP3o2ipP1KOGOINBjiOPyAa+npCl8iRPJRzxarfULWbr6rj
/TYKz3zi5U8Uv/zKw3aYnqwbXQyfmhs1wTjwc2BDdwviZwr4HDwf1hmEccAgbUFmPd+fx7r+jGYx
9NpRc1iFBbom+MYiW5wSFmp5PWaLiaNfqsuP151xbisvbd4E/NvYCIdZylb14E8BNNoitYdVOd69
Es4HZYR9mC2KNZJ5XF787LCpmP7CF/cDNw0ID8g4715on/yoBhEkQaMeBaZjyQyuWDho4RRzcRdS
zoo2ljN61ng/cFWt9FQYHjjkK+lg4BfJKQnAzaDPxTvcDVftr2V54LIxea7wvwlVntZVbMUStt6P
AwQMCiMykCf9n/Lzy9vxZpIjonQRFh0+NFuQSkYUy5qTeEGivDfnB3R61U5GLuGu+kqtQnZxMvAU
zdZiLapXwqR4kAGvFNbdDqyw1r2fI/UwDfXgqJGxVGtliJTORRK6sgJxxdIC530AMCbpPOGAaYSQ
5X9opeO7J1EvLWeO1VN4UPJiY5dUEVsDuOHJH28Lm7666kAGGqzqoTLM/AIkARLfi93Cd918iLA3
tu9sG7tcTOXc4wy+oDhp0tkEkKh9lrGYc2W4lQnocQIthB28+rnOVlA8iCgoB6ojHf8HwMi1FKkg
y5hEeakQNr98Ng+lPs9lzHebPOTfD0ouKxwYn3BBp3uA6pRXNaEseNNaTo0+ImfD/6jLovddWmcA
sFC6GhZtGEr053d3QcPu4gIoLp4sPBUmj0zfsP/8HNQX5rJ46b01+z0X4IzRZAloVJYSqhVyXQAO
JSRuPImjWSmi9qCz87yIZWV+umHgaWl2pRMNHXsLxdhjwaww/G8jCtqxMNIvULlLhzZ28mfidoTF
C0GfDsLM4beY8QvVaYjNk0tiFgnMPNSZ90Dxhmu+0TnAy7zFSb6z+aTH1Gcv6FqIcY9jsgsv833b
Yam7hxQiZqfHCpOucIomAqfW6ebqsfiaN+mKn9DhAic+0eOF9h31D6pc/nDguUP/pTcgJGW9s7nM
mS6k8U2/plIl91DBXFv7UfXf1+nC6jssfjpNibqsOMqJBlzKvsMF89y/sAjFx4FML4rE97vbCZlQ
o6BD0kuxiZeBJcn9tA8yuhJvey1QqMutmpdXFTT/78zWjpbg810lSD05nEN7OBR5v9EqcjHJKJiU
HY6/yCHgQyL5Wfodh0gJG6d1FfBIFn0ehm39WosDYVY7zDMCSMeTTNjMcpsfmEpRGfm6/3JLWD8v
agpXK/u90LM+wkQaIDN4mfE2zvLsWXsq1snPQ5r5IKHEEMwoUPeu1j8vi+QT+ADiZ9CcPhWReD3d
WRbYjVHZ58IGi4TzIR2t7VIFbHHNpAKedbH6KSVfxF3uGNfilX4lq/VcBdTL6qlKmnJHxTaMJCiG
9STgycQCthaRG3LBF8ujuVsbLKGnjC5/8zBB9hU0li3DTlyOPK7Y/3kg3b7oNYUbwlhyUz3RWULb
5grt4VjIdLbCieQfekFJ6ITsBsBNS8Sd2R2+CWclAT/EMkLezcrxrXunjY+4QNdMDlknrb5AvDb+
gqC3gCvVEpDap3LXIW1nAJGSZdgXBcqTjIXk4q8RZCx2EJ9vXWUisRgWugkjJ9GMfAK4+0mwYO0d
RSy6g8bTZSqP9N2e1BTn+hhLP9W/xME6J1tKSVye4puWefYUtGhVwTGpqNweBCpH3De/ZVRONga4
weVR4aTyR/XWP96qB5hZxg7PkYiHGKmk1ocp3DrOdwv7UUSCsZXKPNGuln8XP5GjqK5WplW5Qly2
47VXpdlnOF7HvDD+Lykm6fI+OGjCFdPakqGUYYt3CY4zoV3RCXqL3qZAZRZCXHM/681vek9bkMs2
PPj2wCI3zjXVVLJRSuB9F/FmMz4lYWYbaMOB5VLP73SSrH/de+hYE7VQVP1xy6QuG8ePFFY1N/s0
sy6iYSDxjNh4iO5VyggSXFOoRaa19ARp4jWwhYRQozKzNcwTNXJkQTxT0x80r5JtLtoBgvEHW/vQ
vK8oSy1AC6KeFnk8EMt8oGp9EXtXDBOudBM92nAsVHS6S4bLD5Grwb8VwwgAsyIAmvXLuknkHUXM
m3eXQF/mi4XBR5D2ZoU4u/8VLwocp/jyirJZ8x5ncI33M/x0+3GEOC+XqFVv/GPENVAW2boI0GGQ
H4k7gcH0f8R0tsigpSuocQ13bC0n3BpZO0gLDP3Gwm+19UitkOhjw/5k21xmdBzDj+q/QuHFKE4r
3yulr+LzWr+6LWMuuj3jT7crqYcO4V/V2WS3HeFG5Z1czt/lW/F6f7WX03tFJ1RXW1TwnnccQcWo
kmGI55tE/CohitLaG914U89b+PiUnY+9HD3CWmCGgJxbfXZjWfkxydfxD0n34wN+kx30+4o4Gzvy
4DENhnDHDwH3I9FoNoxuv0hb6H4HBdrPpEeX1nzNjZzUkF1qlLl7/ZM/K45HoBlg/1scPCktwezU
fst70xJbjYSsoPa8YO5x4jX0Ai+yRKD1onr0xC4dWlz3htFHQL7z/ea/P9/IGb060VHwFcn57+gg
zlDD2bzHxb/rb1vVTog8XcQpeXN0H3Kg+BMnnQ3R2tj8C7Lr2e+tCgpb6jYsccTIzWPm9OKAIhs+
sPfZGS6stKEi035Kxp/oaYlWgba0jnPohJD7fBgsRbKi5LoZ9mbFx/r3pzwSGnsxzjzwkQlQM8IE
FEnmV6OZWIqu4vqKNgeoJr3xP9jKSmE33oVBGVFQIb0K7UmL1HNTbonROjjPa750qSmiZkJ9rcVZ
MxUM5N+Bp0eWtAo+W85Dl89oaKwprnmxqfJ9xIZYFEwsgM0GPH+1xbqhbIhIWBw8OU19Aa4IYvto
Alikwa729MGLge91sFNS/i9M7KoEG2Sd7YpvwyWdOx2OS4BqkTrld3Rs+L11GhmsE2PI1DnY8bDy
eNAHtvsMGNQC3Ed0nUvyHVV+xutORsUDvdIO4BPLsoVamEbHR9g11MkCY9gcRVfojxawAgnwk/0h
ZcPvMrui22IKU8pcaLjlDj3nNtFUz+PvdxaN51SDZsDpID/s4VzHlfaiFJFLYSzGuy0ldwD1Uz7w
qJqf4BxyLF/4i9773azhnNhs15gvDbIsMgic9REAnH46dzkBvnwHSb0a7lRQtovj5oSFkwRXRU6U
c0DPdTCPDXfKOCeYkS93zWR1XZWh2hu5GXtXcnaYPVNQwkyvfUz73xrjJfgEEYcOkf2AZkzVsjxI
/GREJTKupWik0LxgAEKBZV3TAGJ4IYuOGi+Vo/2pmdCDqQRkWKpdWop+ULZO6ZScNMp8l43ASnX2
pcPqH0pmr2zOh421vjhRzrvY46vGi5mrdNt9glwPrkEhL54/BIWLgDIEHXP6SCLZt9LUxIi6kUMz
gaYqTOW1AahvOWWxkL8Y22dm7cO8R7EPywMSxSFSCZR0tnVlir07CgddxE9v0ANq7sTpvIp3660Y
Vz8EpCP77oU/vwLn7K2A3ngBiTE8m2F2EnsBftnYHlceidkhHN49i6RsdMFOhCwTW7feY//meC66
XOCkGCZO2htsDfqeO7Z+tOxl1ZwnsltLXKlWvUkfYw/mdmcLmEUukYJxez/Q1V8WyumwbEcMiqRS
tkCvXvqv2h7WY8O1Jam2G+2gMR3EIuUUrOy1iTYXsDt2J8sIBOUNIb283XCIP4gmogJc4/ucK62/
i4jMLfcOktgjPwlvVcKEtXa2DB0gjIVVl87Pp1iITlzsrJf3VQQ2j9dFZbCcGZTagVxnDJA73+GQ
nyjcdy7yavmm6fyIX/txeJEPYS7z1PhV8LOw9AMWexVEtHS/+8qPrGHa9xiUWbI/itD7bZFzJ87p
r/M34KB7vKmASsr8mrFv4mBiZpNgzqarSEZIGedOtZ8wY8cqguwxXOjTjjOVHXj8GPwKS2wdQJPY
mSQQW7ukDOJOh0ZvpEApA43hjZN0jUn3J3Jg1n9DR8T+14eBEEN+0iYFWZQT+Ncc0AzfOP+Udgzy
fxh905tSMTST81HypW4vRi1GOSCDWpYBksrqmLrzk5ZNqRh5XFtdJPMaewRF8Z6mM2+iq+6Qa/i6
EHSxKwm5902oFNJ3j1ddaezy06mqy6FoIUZnby6pO8YomV26PcEv2RT2qhXOkQ67v8Gtc4qHLYfG
iiE9C+LZauwO2n+tiCfs86IfbOXFiC0xbyrMKDQ/qY3Tmv8S+ZpOHAKxZ5bQoYT2iBcBJCS+n25n
1qLtWqxFCOmxLo5Qw/b69K3DammlVkmMeNlH31Z3yQmBGvR1A4bh+0fscYWISdTkRKTi+7EvycKt
zs/O254ncA7JhsKK3MX4oxT8TRrVjjnCdvsLJL5ZqcqGy1uUsGInmh5mYEUjas1eifkNMv1LhKYp
c9+vRXF4iA9vqsSTyHC1Jljak1kqliwUPW+83FGUhR0IeHRea2FTA0dk0SvCEteOZ5E1J1dfkPKs
BGTqSY9uVmHVcDiUmyyQMNHBGItaqy/HHkTQ0LiNSQjL4F5nYyC7j4A7vDyYHCwmEvT0VoFZOcUp
1p0Bbg0+DcifI/nug2kYBTycTTj1+lsh5Ol76myblVbfj5NZM1XOJyz4LDF4ALJzt7O9Rg9wpQLa
E1YMZ9SlqQsTSI5ln1ev1WMx09yH3XQL3OzF/+LKHSCYm+b0B4c5sSfdo9coFgNPNNAv8wM0qK+/
+ZmHB82+qDdWODhLAtTlr0MlRCkw4Kn0DXmMLowB9YZ5Wzo4fwT2XzHNV1Lv/ifm5oiJBUEB7sSg
JVTumEgtGD/2ifhoT5Wvb6LOOjgY/jaQmLidsQ24I7gKkSg5b7AarttDlSLIxrnP9QjXMavxk4iw
+o7wHO5/2lX+vI8BPLtYeavqmll0cZS/OBSIEaZ1ydgfGwmNy3JoT8hUsCNLyHC+095l8lhq99q/
y6NM91iPmsBbLxSHI8+w8c0J9r+a7NOkYsmLKEteOTI1+PsaYJ5KUMWnfIzPO2G0d/QQn4JkH/oh
uk1rkN+BttzsBdgW6fbCzeifHiLTyKjiRmHc0Ts8RpjlVp6i0eD4Rz56xonhOCdeHoxNowMv77Pz
QL79wE9YcAIgQhOfFPQioBqi5eaD/xjDyomvwktwiTto4cUCn1yKdOPyILCmj6xtZRaS6ojUHeB7
dnGep+jXrqLrnRKwTDDHpO1qg01rBMakytznsEC+EFiuzOwPTpN01a1l/fdMmypyFqXVcybNB+Lq
yYX6MSdoFj5GNlsucTvMzbKcUD6UuxKq9uRFPyTtfcre4VxYZrBCbyofEKf6hFchrxrhPuhnJpUH
ztgpbjkbj0ZDMUG4XFFb5CRkBQSBpLovvOhZwN0ipBUsals8KSry7DBo0afBL+xCgYdaypodSgXG
nK+unAS4VQqhi1kzG425LgGMt2AIVqA7dmakjc/aGFiMkvlVv91u0u2Elt8F+lnATwXIMhymdBel
d889s4kC5UjUxQDa6nr5S+uKRzimrPVhXMiIVbq+MR1gGjs+xAU+C4VGob6uEGq+7PXFONb8dLBa
Y7j6CBuR62dPcWex4qcXjrTxAiFV3L6xBzlLHDV24yKjgB9Pe/9Ci7LQEgv4zP0Q1nZQQpkQZr8N
G/sfKJZATbEhdowWS/jjT0dN10aGDC8drssGU9ODFLhlDSkC4oKU1AjBdU5MPlPb9GOiINS8gYKk
dGcGD+iU0hv7X61X3TMA5aKQMqcxzVCwJt8T/EtmNcyalcxYqQFTx8vDbCxrNXPTget6PpMSbOYP
RBSMJ692rLQsRW2xYIO7qgXZnwnYi1S7Srcws3rOAyMy/GsK9wXN1WGuxlZ8r/cTsIJfQSR8Xuv/
SUN32CZQ8s2YiWYLnExsv/l54xbUGKzBsOfFD9DeWaMaTBea/+8QCpJEbuDvV7mSBEAeN1qUoMmc
fI8CCSiaFEzJ3E5PzU06hyiqKjCk4KIRh8ZRWAsRElZNX/BgoUQiwmgC/W0CXLoVTsIID6vAGllL
p26FysEjnFiJQvilmGSFRosUg4K2TPf+3l6uGl6Fy1dciJoM7x8WfP1eK3n8JGrHQbFkOKEggGjV
XHyVmbP9DghhC4QCJVbVAOU8wbePeLD5iMFCfX4mljHAZbahcJLC3zsobzZ0aEGTHLa7hYIPwQFS
ftNlsdDLlTpmiqQ2J0xAfJrx2H1TLOaoHNc62LQ6zSzpKWzrxxSbR9sXlOb4IYVmdww+Lg2jbusF
dQHFCINSjkEnyuD8MPXvjS7uDlbtlAMORxtFQzUfdLoRX6xPpHdSswbncxIZQodbBLBRx3nErXUZ
Vq76DOm+g/L0eiXKOx7sU0UgLbmAlwC9KlQS5k7EmqMUz4fIeW345QLuEHHuH4HVu6F5Z9qnzDTC
g3pW1tpwSY9Jsc9/qo140U0za5i7baO+KzJOltectdnuqGh4KbFOPF4VrRhahJTstprllf8NGbA9
5M6BjEw3lB8OeTJXx+lWtSt29t/XNspP2MAXJaZjwoG82mcibPpqi16wYrL1rmbQDU2Ni2m9o9aj
VkOEd8thnpOHNT+9ury/zl8tdXtBh1Vxh+KK53NUkOs2XU0DcVnmZwifgUFLKnrYl/Lw+fyiTDDh
Iu2udN/uFktRJGNPT/7rHD21PxS9bjvkkhRchYt6kXZ+CNy49UsMubp3fAwpkChdAK2nCw0c4Y67
tu0Evxgnor2xvrB8SxOhVo9NnGxb8LFxTksukt0ZrHMQnD1TPpgM5felgQWGFM9U48ICZSbn7PjU
inpDHL6qgBM4JgFtZjYK2r6sZk8wiT6OcIDDwz58TxIH2saI5g31NKCNJ6B70/iBEsxHC0NtFuc2
JHub4PNt1qzn6PduAydbfJ5ql0hllJy29PtF1TmAnGUCBJh0bdiCItYtrBdxcjI3LN2IgwUEQlJM
aaXpmaPvZbA+dP/XI6q7dYbvY5sgsOS3IryjVzYhizaN2YidxZdZECZ/MCM11RvlTRf8NcUojVGc
hBh6jAhRP1J+kH1kc44ENhK/X8I5bX+m19ZQay3iws6H1eKyjtGz6qFWnhZl9nWtPXvVq2/R18pd
iQZQmBijI0I9o87LvEJphsIgUJykAC9KVNxoOGTvNVOvIG1jSwzS3688Yct+0+nCwUBlLtPS49D2
7plBrQ1nKDC/2B+E3iUEL1D5YDCto3ZQ0Ne0RLyNHfg3DJT6icrBvwGEi8VxvaOrQLjMG7U8P1Xz
qc3HWWbTE4nKoLYnkUVC4n/vT9zr+47TKdMyd7crU32EsROgvVSAbxEqTAjn2d525CHhEPDqT0Ug
5FFM29sIUx6Reb4PDVsbB6h8p/f1LAnIuU9FA2m8w4XM7GPFZuMedh16vQImlRlh//XTdiw98rDa
X/bg4AoluqmCJCOfENoWTOdpWwxPxyZLK3IK2wZ3lG+MpRGpdM2feBqhFoxXjDqeXb8uOcp/kVBj
M39kD6Th8weUsVQoNNKK5xEWYL/+hrPVRtxuVO2XxSBJtmoH0qsxbV8ywhf0r3oSr1cra0MEI/Xl
B7Nv1Zd67DV+ngYmn6tQkHfDkfUMYBuiR6DCdoEX+TAuMcVQWhFcva99bU+bFfoxA2xcEkYGFETe
nRTKf4BCiaS8vdUiij0y7YVvZIekFDqXJtFoXcStpEL5Rs0dHgkZQbwrjFZFvdw5z985sl8porkG
cIBL3f4J2kLtYBNcTi6PBNaHwiRiyeSOeS9Z+ndDzUTcKFjCsdWXtWv1pBRQd8JlY4W0WTtNIhz7
dI0t3JDwmip4J76xibHwP2NQnF1U4zcZ89LpY6kN1D1Z3a+ZDH/j9brrsWOK/7MOXtY/xuLRG54j
w3Vri6ZMzvR74+jRlqpdPiphds7INBBOhKU7BKBtb54KJHvZnKMbrwlVkaSKdiLJ/JOKJT15VODE
iQtfgVHVjeDRmw0cjK7HOZCX/eQMBOb+MTfBdgStFeMU83pA6KasLGwI5a3TRjhq/zxQ5eFkgMz3
cFMQzcKnUEsSC7+Hk/l/E8yj6tDLFn3kCDa9s+i4L6a3953RfPDrH7D7pccxnb3WKvLhyj4WBdF0
Z7H/G6T9+gSwWSwNdqZ0zwgyfyd5i2+s+Jt1FhrLmE+sFA4a8oQW9rXaSUTOUEVWOW1VlNwQe7ae
/7/1qkwhP9p3x4kWfqjO6D9CvCrnQx3izTs8QRfBHwEwckYaIOJlmzkUYS4JOYmhxEP4cNQZFZ0B
BNkaW6GpHYtOJkc5v00R4LL1fKVxfny3YWPKb/0v+mfaPBnaiFTEMRhf95an5JEyER0P30WOYBlC
pbSqAkz9IQqNkeJmrGxm+jSAK2DydiTWLQmJdqmLHS1Fwoydw27vO4UpLjsn13sUORgpBdns0xdu
PYP9BoRQ+0CW0lNogK9WZ3MfPCh3b2Uw1vr6TIYolBl6zm5wc/y1RPo26rH/UnruklXo/08glGRq
ygUZ9GMDfJfW45ZNr8f7XkzpknjozNw3dnFSXXRaxyIOe1UAsh8XaSefT1xdb7ixvxUbZX2XQ6WB
bQxHRWV/K/RqlOoo+ukqkrP0pC4mhPthjMdlLWew01zR2gNSwfhDg1NL8cSW35AS14noo50VkP7k
zugIqqUj8FxNthzXPeZEo6R3tPknaSJZQ2nplZ4dfdFp4LDZ2iTJPFMV/2Q1COmVBNMAkKrk0JfE
Pk80xFwaQpxBrEXpRs2aHp98b0fpqDFZVmdGTwbvauaXlgJ5r5N4OwI5TT43py+rN269WaFe+LAt
PPcr0O/Yg7ufCfdiGUM1rvx7zAwqh7OG19Jtsx0Mf/S/wtEnK6mv/QDyZqpvj0XH/T9Z5tJPLDOC
1bnrzzAoGO0ho7eyZWyT0cvdzsMbunaeDeJKEUslObxx8/AwRu9mcanB3N4p17/lZck9px9zzj9v
yKuHi+e0FJUmF2BXntdjFaKhqKL3hfqClI237t4U7rtwobEsLMni7Orfz5VVb0XVVQ3tgppLWNv+
PKIqWgFg4lTwhS79BtRrH8s02JMFS7QOJ05kvoEP1FLdCsIwOI2ozwLi+qLz+eSv2iGvXL9vwdmQ
MGmaoKw1N4aQamZc0kQPfoVnNwVe1lmeW7EQ4TmDFpiY3ln8AF/9t1fuE2/66ywcmIqLVtnrKYaq
Wxp9X5CJ98haf+pJ5Mo7QYEs5jhTtRp5NhEnOrCjevCMLQogqjELpQNC3fMrkkrN8pooUmre1fkS
XCctIRh6R0sU9iq66xVKoJ/VuAUFy+p0TwFe00fVoTv2BZHTVO3vMF01sbhTwQeb8vI6pJkmxKvc
VvFyuVj4uePvU4z7CIEiP5mH+NzyO0lpmYTmyb3QDxAjVjGGN27sWSu30Qwdb6WfF2WKqGT0G1bZ
8HZ6z8fGS28rPN/773+c9w+cd2PPlbnm0c2YZ2ZBJ3cf2g7tEpNN4n5DVZgTFPwRIJAYPd1xcO6a
12smlX6Cr9GMs1hLrJ9SM9/qn9ymUUuCA0LeguBt0jGoN9Uo/d1L1KpBmBN8zihpP42KoUGcdwWR
rX1OWOK2lnJqqEL4aKDg9HL4GQhpuozjFZ0JdBGN2HIf4KwRIdct1hLAX17cFxBHe3pwjuhKE/W5
TdOhRUxcpTwLEAqiQKMNR9Us62NONfXhx4gEgBGdHYy9ckt25fwB1A+7nydp7y5X6txY07tpPjFe
ob15nJkHWNztz4muExn0tIwKWTpwyAVHmOr0MUi2/77fywD4MdUGOSgjt1ZtyFnh/j/E1I9jPE9U
Afmx6ocZRrha54ExFeOOjshHNnAEK7g0wbWWhfJnvT8VrpjY/FF9Gjppw8O48JbvAPTYYQzPpkaZ
NkBduPq+vZFWB1wezZcZHQSFhB9XBRzN9c2fWjpm0djCGkMEoa3od8ceFmEhJIqnKCbUOI3MpTHZ
kjQ8X2K5W0mBHv+CGu6j29FFkqEQdT4sKoyjhuBbUeyby6Y81hokml/XRnSttKAhSXNeNSGULjUM
EGp0t8Mopw8MHJ22yv0wxbOz6mOfvpJACrS3sT0vyNipXBdlelvuoPERuCnhcyIEFIxvrIdQI0Y8
0HmRO/w8emSnAGYOYosByQw9TnPMpsnxiNeIj7bXOCDpNA971H58VG2OxNR1IC/jmGZT6MpsPxZ4
LrJmhO5O4BPXclmMRz6TGzONrNBPYg61bCaiCgT6mv3QOfBXrZxBpnKssAVZgZDVU5xl0hws1INe
Nd5EpVDqte6kfWNFrWS5LCkHizUw8Ibyly0vesGD5iREkLcEEM039KdwCzWUuIQTV1CpomVDWtEw
jIe03wDbYDjJ/UKXw0mGRBvK4mHCo4YtbqUvq7GGhbJS7HuvcBUSXaHpnzLG36ibHD+adk/Hlnpc
FtzI8OprQsBSqDHA1PcyWX6GY385ZhNAhSEmZZiAOwmbDhTCbTLXRvAjyCGy91ZE+L/77QcRq/P5
vTo0/9mqy4bNYQZ4VTDbEL6UDr8xZTdxkCBV0Xd6+jl/eln5lHLXEgXGWmRalz4yoRrKh4/cDLVu
57yOc/TujkGFaIzp26U2/jsocj4dBZrMAj+0Uu35sscuF/hjPBbE/hKh39xIr4OBplAWE+FDN59R
iapViS2wR+x28MiZrWiKUddmZp1stFPTxx/7XtX0z1dCxBT+voLOzcCziCsGY6zgahnKbUjLTeTh
uB6qJAuL0PPtaM7KKPSdpPa3XNFGGOIMi2z8YJuCK0s/LEqV1I3V+ycfbO1l5EE67uY5rTfvRNwE
TfUOJzqBVroFTPOLKfLo8GPBj7t48jH6mYqSA4fXKejbWSLsw8pSTRhi2djbV3Zll4neKXoLjxAO
jg+nqYgklDYAbke7pFH7TBU7tQyxd13vcxEDM737CZecfYq9npiYcWfhnGL6LVaMnufMLUUFKDKQ
iFhEwc3/8kDAECxT0p5DgdIbxyY/z7QSio99j5sQgCBKWE22BamwsGn8qyU7Z50viuVDC1jN8BaH
I2f9vPlfL3dKFnqLO3IjM1bgoz/CYY+YTSaOr3BgZ5lepVlRYuAm92fXfNKB1rDadwDNP/EhRtLH
LLIWuHf+G31FxC+qAI/Aoxb8a7l0ctZ83mAaYnjCIgGPCAxTIbUS9VbOxLlhEzEB5DJQ0jhP3MjV
rsa6Gcg/APvxx7O+ueK8+aiaPp0BNSejeqRXDZGl8SjfRqa2Al88hkKtO/mtztjCD+iG/asdXxLy
HtXO/rkJhyNPdg99GzKszcjG1M8626Hix8VssYvb8kQnAZBJWwvwNqtpWo1jjSolXaa2lxl/IkAl
4nt9mQKsgP6eyktlBNBhbRyDPCDNsaso1RNW6m3pTCaVUEscijIv5ncZm/hbH06D2XOk3xbi0pVj
5w4uT1t7+XH9ypLsz3xLkLSAHcBLQrmohOB18EnIe7oRrEjXN4IDaU+f/ec9JUiTuxA48dEdv2Gl
C05R5DJpoUi1LQ2Qz+SaylL8f/rcx17fZw2m/cuc61ddXXxiMPn9oooHZXEEBAZ+eQzzKPD1+ZjL
aSI0ZKkV1Wcpow64Z8ZLSBUhdtfdMoZ7DnwFgr5mrK3iIl16SKgjUHPeZ2+Bub+9r6cUkWXYE31b
9td1fRR3oDv3RGoUEQBgJMkOIzwSrgNglCJJQ5z7D1RWtlvQxjWJ5x56M7BqiDudRZLVVfrsZA7J
aoXm4JHJ6sjcqbAL/iWaVoOBiYraqSfGPYuWjVjMOqbVXAJU4jNfZxoUk2J4kDzpebdZ4d3GzhZc
rZBkOp6rxyJ4nBvTKWP20/861ani4NxgK3tZRHMv61fjHW/gplpKBGDNGaNbSFjX1gmU2g78DCnB
3FJZaxDagL627rd5pRTlcgFYZ6DOmQD+Un+Xd8D4MNL9pdSb0LA4KXVozdr4V8z/vgRv6ucOU+s4
WQt5mIeg8oJiy3z4FF/MSW12hhMAzXbUFOejhCYyAZJjPJ93SzjbylJm1MKd9j1YAtVvLXDY5WGc
4Zzzbl2wqN9lCCETbINnCzxqP/1dXjGNHK8sGA3vRoxGjU9CCKbxP5oDP8TTZCeqyUj19Q6oST2W
IMktkWxI7T0Fvi6cnrYHbxrJ4esiTJFCcJNWVA8MNdt3IRbygbX+kEjv5Zkf5NoaFOtAUZpt0xql
XV3UuTinJtbpEPJQL1xlr7hUERw4BPTSvpfeha5dl7dzcvw4Swbz0HBOf3/A8iAJbULTHMfncpia
wElY2sjn5yYbRMaoSpbEwAnOty5rRMXKzfclZfiAOA0qvK3ty8oqB+KAhIeF1fsDmhhkr+6zf9UV
oLGCAtd9/c2WiuJN8XWjKtOaM5cm8xVkx4SyEaKeTWQvcta+Uwx5ts2oMtlKysoKVhsnaw6oirCa
iMxp9tB5BV5XX1bzAiHrAhR7deGrQvmfR0tHi1oFX/XU7iYvhDh4v/Vo5C4bo2FkA2Ev4nbHoMqm
/WWabgraCSAmeW5ycBU1G2YA7FnXmGhyUXMAt1VzPN6XBhUWzlXHVlbWFhztjCPlUXJGuM2ake5F
WfDO5D/supYNh90tJOpIZRMB7LXJEuDPf9IJGhgoDJavqSBgJ12enQBtf91pyMPEBVjx1ON4Ayy2
91bd6LvPk1twiPqybx1YJwvf0FKdy+lhXfLOKU6WsdDQn7hQcJsmN3dsD2Vzn0xLHVr1dJeeXNTQ
6R16Rrr3LK1HfjabG/kg9GqfC6s3V1Hq4hacft9sV2W14VDFCLRQR4NNlfOvh17+wtw9Pk5mpjZl
lO4N4jELKIoMSrGkH+oalUMvuYqvpTTaJ/soo+DN523XlD0OAjkDyO89knasOzKk+S80mvG2rmvR
NgCywvG6uQXQJf/q8dIZ92I8vPtNolq/GE2xMmUOppWSjN0iK0yD7JikpYU5z0CC8l5vPS4Px58P
n6Z2CWXbd67pKW77XgIBMm7q318kjyW3DvdU+TqSCOoCVs6VzkD5NilKxJG84OGDpu3pGCBaUz3q
Xfn/MhhejuE9T83JhxIEi0776UUL87GrIuHShGo181EXO35i4aE+nzuxXedQgKxzVPutUqIosTB9
VYxouShHE5LNZQiBKIbYO7GyYFl/fIl3vydGP8rU3NOT17Uu5BbnMoDefk+OzjogCs8qaN5WiPJD
b+4d8bhd17tkJprs+xZ4vP+8tDRypJ13VHjjCYZx8AHbkvOyPNcS6AFOqx5Dr7L4U7CDeFf/8Xz+
pLfZQeg+If1M3STK7EgG9b2VdqOUFyx09sMsWdTN/VRECDxlM9RoLUG14FACpQqaqL/kFOnI5VRB
uUp5mwXozmLxytTQ21AnDf2nra0G3nvh59MP9iSe4x1NNlxcbV8UqCozEPovLxqKcDOyBi+xnLbe
hNvymmAWwE1qSzN2EoPJ0WMij8Rq8IhoeN6YmWQQbJ3FKXVN3fg20u5Cyc0cyUoEvw7JBVDIMisX
leWmnGd/lz2iGpewYl9sg2GADsZhpg0mo+PhalG1RJb9b/pBJOQG+dCeshihOneCXXysPx0bMf85
cnwhb1MeSallpdOsFhSWS/w+3YnRZtUPOzfDawBdwjHij7Ht8dsoC7aPx4hKEyUVvnEob8+ic7Vz
FSSfpFmDhd4O3P0OUU2ZJ5yOmynOde18q7V0HmB01SR6B43Cd1lPF8vZaz8KX3JwZT2NK5+0hHSY
yKLSdh8Kis9HVuBfi8KzSXyzVcaJ07Fg8zYVXzj5EcC+35dWbyyNnIBj3DxkSFNY81o/oIxfxHIJ
ATF799MLL0x9d9/r1HeyoiSOKmAXazok2c+fHwUa3dtNwq9nzZhAI14uozBkwMuEpijMW56YT8Es
W9WkcKEeC1i9Ps1w9ipKlAoCzZxlmsre2a9nkMGVNruPN/IQBS+pKlUH0Az+EjEnd4YpjJmeekYV
1JrrcFi7gyouAocs1RFs79cbyv8g8vX8B4lfGDUdoKtV6La4ilWsh6IaW00+8DghOF5EnQ4EVTnS
yOawc/11VX+BtjWItfawA/Ug0wQ1oU1SEdzFLdjZpoMe3+1LOPCfL6jmloj876bObFXWoH4Iigrl
PO3awfOMPBasIXZKwlmAUyIDf2yJICMswzQXiojVdg9y4+jRqvYyNJumuFsXMP3WhUJ8moT9DjrJ
6/VAYCHavhvdmZ8ABV8jUUpwy3AxMH2amKMVyVBK9QpFxKmgLLd10SY1n6c6dqMlTB3o8i7w5cbs
EaVxdcxjUFCr/yBK9+fQBjWva3aaFhiiY2exFxV3SXwQfGTtPRQqvrzJEWpFRqG6o1WJEhttl64d
cB6vKQ5yUS0FRAwg0KVudDXd5uEThHL50fCr8fWwpiWzX6/dqSVs7yDEoW9uOFcc6u6jCchprjvR
kVrEdfmmZEjwHUReO4gMAH4i/9qdAa6gmMaf257L4uj/2JJe8VaHRknJYDSOrMY2M100hernJImc
pxlSfEG9R9KTGecV1Je0CTS44zz2NfRsdRbdcgPZ1bQJ9EueVg1MV3uwRuGUCU1zGWmd11p58n7C
y1qhc8qPCw137+SxvC7xkHfhcVRS3bb1RKmSnykrvrFvsNHqLnXvNMGVhssOC0JPL+o6Y0ak88IK
7qLHUgoQ0c38THbnjWCNXFPoGjnmUFchPUG+f4jJZkLGqOisPziBxb8iZx+LKtR68Jb0nCmS7Nev
k1rpEBoqBTKalQtKoMml610nAtIpXmX1TkknurgkWgoqvO1stwj29dQwptc9B/6tGD432Rv1u1z4
ZUgjtu6hihgvKOLi3Z+9w+YwW1h5d/d2xdGX+2Iailo73pGB2bSXl4FqJ+4eB7n600NadETzxPtO
GvIyx3l9o3A3t6TrdjKTawUvecDUAPiar/t6ayraig7vW1AstXes9sKxGf4iViAZnDC0AEdJVReu
E1fmjCUqc0dpsM53jCAaqMR5uk9Klw/2oETKmfKvxAfsXjFu+RjTGdtadcTGHAk4S+ZQw2BehpjZ
dK9sUsSPakdXh76NSDzi61nAMoNhsuFayEiduvrgCvgME6waIEcqMo7qLrtQpEKu6jZq6OO5KOMN
vsTNC2coxT7GO20vPmxqKnD8DXzOVD0EjbLMd1IL2/7OsuhJEkQNxtvbQaFgO4z4CpViw94EFSR2
bRmam/TBlZVlFWg0gVlhEzcTYvi09usg/bxDi4ccMV9SJTb+o+cy/UH5T6KMjn8+S3qmyjMsM9W6
9j3UOJ9qXHCQyAiowsZkPUzgmC/Yg2+wIRoUX3XEwFPMpJmU2B5gTSgGLOQE1WgsQ64kkZivZbAl
k93GUfQNqv2ysSnUrUGw5FnSvwt4ldGaKPpYLb0E5B4OqEw+69mZDR5WuXADz+4OipA23tCNY2pq
zPQ1KVOrc+EylItiSDXz9TFG51odX/snainm82RfQn4WYvX+RqsOdl7Pf+g0JLwe7aunYxqDQblX
nrAh3T9/XoMvzBxQzKSvfZ33OxhraTodNw6MigeUUTmnI046v8d+esgH8pzCEO2MjjBX+QEk+8/m
jhuGVsv47uIq6tyun4rHbxnmK6REuMmGhlNXdOscAri9daa83Gq6zAiXRpj5rx60YtIdbsA1wEAu
+uryXzAgyJOVWp8LcqkDVuh7qP94YA99aRcdrX27GTtw7/3LtFbkczSir7mn2mrOforxjLKCwPgb
gkidICC8ZSLmsNmDGUzecOGAJPW3pkLR3XD+QKM9NuycZ8OEmPPKg3zhKtcW17B9OS5/vcjr4gF4
ofYqO2jSZucMCyEah88NJk2ihsg2Xv02FD2SmUJ6QF3FNgZ0by8uC7VMS+LhltIv4/nkC7yCpxR4
66o5LbHIudj9FaRelopppZQMId+HjsyW7Thhk5NlewZjfyX1YQYTHPdseXNM0tx6o0HUUq5GIBaq
FRDXKDnCa0GIbTQtpupNE1BePoGQxxbeetwaNhAqLit4rqr4TaQPr8COM0uQEA1eUko50v+tBEEF
aKqnjRHKRZ85OPVqP+1wO9gjS+8tsX9t7IR7eiydsdhr1D7jIypBaSmUKpQ2O/KNrAmnbu5CHGCE
+twa9I5L6neyC+H6K1DnxIYqZ8/RmiUPi5JMOFdWooyf1hLFRUUK/g9w5JRNyQwz7MNDj+aRR4q0
/d0SzIDgUJyOCITQqgxKQjTRI36i8ROpVuC5Gty/Cyws1f8BKoL20nvCQSCAZYZXAqujSY0cPtkV
HEM3GW2IBJClAWo9SHhczAROU+dzdkuCb09qolExYpZBi+zoxc13qiOHJ2qyS0bEoUo+CT44L1fU
0/OBntrz8OsQJhjngpX7B6Wu4DgAcmuOQeuU4s0izgpKCx2Wa+/dyCyaV0tj/UrTMvMc2PTunbxx
UyhGlZqiBFmlx8nAxFhl2KKCcUlDa8ys/XYmquloVF7IhoAQrv80RBvP0VXF/LY9EQENERZ7a/IB
GYpTbaPN2vKIOqDlfSZGaaUGXReEmKQrHNIyg+inAMGTu/5OWkv3KlSiQYrpZwz/GinQ9tqoMwsq
STPYf2Br3ZoRa7Fc7nHbPIRr3uVA120ppawAZwTta4a0WfeXutLSDhyKc8Xyvv93Yf/c84biqSaQ
nvDifPdwZy59bF7VCbQWSREH7W/hFBaGkHMzeup5m5fznllf8rCsDqnKbQJyRKi/UuenbJRTfDKe
eWviEaGuoTvfCMApAR1pz7k5zM+nZxnKFKIqY2ei1AcwSDHjk0Apgtl7qTG6hvMUYGb9Xm3Qy+kV
GbNEcwbsE5zzyYwS8PhUlEF0SXGOjcrSSKrkSA1rUsM15KFJBI0rJ7FNVXvMZBjnhaobH5u5qPhT
IK9oCZGdRyQ8Ec3d2l1W5xc0YrXpWRQt/5JslFNYNgCLuNkOtOxhhlpaSNOu/Szd56BYYqw8HUGz
uZGxjAvU5an1pBT/GvR4BsWcZMHxSZlEVMecp4RZELgaUchpiXjIMunsl4OOfsGnRNbiSoH9dxgy
1dQZPYpERC3R3Gxkvwx9dFvnmj+x7tWrYQkFaMSQgjvIKJ5vj5+H1zoayRIHHk6+3RdeY3RT1Tbw
tPL5WMdbnLpk14ar1ZnvwFW7Vgz5QZtEkq8qIxJlNcYU2NLxtZuS61+92ztwJyd22CqwQKsCU9LQ
E79t544D4Jyn676UwTtwnP5xEypqBXuTOZGokxbcMGlwR0NC8nsKIDAImI9rF4731/2osIT8zR7j
x6+3n5ZQs5gBHrfYRQBfuyXS/LR2ombskFYsFTb0AptYJGFSTRbttlZRMyevEJ/SzMEriSx9U/t8
BgWLM4gb7Z3mn22YLaMEO7HfsTxF4rWSr6up73/VpXwNmJXYxhEst3UmHbwUMa5+AJCsv4rJqGvh
9iA0ejA9D6jwEL8oIPCkOi/6zd2UatrEb0Pl8viNuOw8KFR+Xb9/1viIMkfVZVJVo90vq06vVIBW
rc4QK148w0I+gRD9FA9OTrz0e75VARb7o1HMFcFJPS8tlcasuwMRsp3HhJOqkQ5rD8yUK7dryBC1
SPp9yIiEU3sSNsemUTv/Zg1FAFn7H3HSXXawFs1qD+NvPTXNTmEw3l49RcH3VV6sH8h906/EoX3y
oqu4YNa8Khcg/RwaOVzazB0G7y4xwYnqZGwt+zv8dNx0jjY6XNUQzm9HX2D3RQdcoVpuVSn9gS2Y
PZXpsrmQHfMxAhyA6+GTzGlmUqDJOdCcOcYVGJQ6+D3LkeWLX0tu36+bKru7qylhaUkxIEMqP6wR
yj2eIBgpxAJ4lbD4TXyIY5sRkDtPcgUpB6i5kaCxze7B2zEuFrXJqGhoAfhx+dCXUvs8jLFp9z1o
SWjBEMWCwLt2qc+vvjKwT3DA4WRvaJrnsrVF2Fekg8bNfmeMcB3iVstsGM/8KLd8Ykfw66ROG4AI
fqszeiIP8630aGupNAfqwnTB5vrdYq8bnuxLMBw9bp7+HsrS3ZjPHBo9i5hSxsL/i4NS0MDyIbL2
yfTdrQpqp4KL6CZ1+Ru43V6VuFuF3Ump2JwUc+4EaQCaCRqpIlhUmtszQU1tsSpNlJDbCx1IQvoo
RxaXEfBYiN3erF8zh9jO4p2pRH49ONg9QOOukW+oUQBLRs8MEsVpxNtg84WUR91U1IfclYV/oGFa
pJAWoJCzvVx43hSj/v7omvGTSEGlt5llZifBQsRApp1WZeS7Sp9LB4BeiAfP2QFxjjVYv06qm9KA
/PqyIiQ/TwgYOWrggkBYmwjL/k3pl2HR9QzNAr2wzK/SF8pixCu4pmAHnfNGr4AoGunWZUHjaq81
FQXogZGzEBQ69j3qmy37aXkyklfSIf1xJ/17LRE6SWB/8V/Yd9+SsqvTXpHLscFKoOUtyaYNsyKk
ujm1Vv0TUyRUmbaTcKYbhguOttW8gOFJqchcqrHr64/bPzmKeO9Ta4IQuge04nFx8BxoPRsv1PgW
IG15T3CFy0ZziNyoO9X1xWc1k4TFj2EnabJ0p+CM6gLlwdICgNtNuYRSQE2OVLLIyU0LrZqnRCiz
hym1fjW6lPs91245EICWV7Yh009nbn68KkLBMJ2mOBJfVgf16FWcI3+a2fPNZ+upNDLzswJEY6/w
zS8juV4By1BXv8MLJ012tzBiq9imA8cwZvjEw6C9Wr7Avum7AHiPLyIy7UeHQ7o7HEU/8ldw8bGm
OGnqsTYz7mmj9WJFoN6TqogW+66GLqUKj7htgG6hmmJXOhfNZ5hS/Gmks5BJLBpz8YNzodQmRE++
c5+dO3IoNQl8PW7YVO8qA480CBW/2HzAuYqgWyvhzbOAPm3Qv2GRzm6vOkVrw4mBoQ0oYi3tnmlB
w7cNLPnECNkRzMA3FRkm6d14U3lrumV5Sk9m25NPkkwqwRmnliFdRYmEs9oU+GOdjmEz7XhZBsE9
WqqTGS3smB7cshRaPDl3zxI04TD68a3egdZj61wCz6ypIpaIc+lOVg0H8W8rD+IHZftCaymLh+Gu
5ykLjyhBdB97o9GP4Pn2vlYgjJjuvyVUnnLu//HdT8o+pa65ikO8wZwJZFUxoZ5NnygnHpTlyLkv
uVeUYrfwkqfTjngd40ASO4jPztGY40DbbqfkL8MfvWUt4sLeFqmNqkNzbKl5AriZIFBil76OOVqe
HgRAtW//foSUYTEuG3doZMBohswSIatWpacCqzQz9h/yqrMKVBIyAOp36yI0x3FtBDQxaWn3nR1f
62XcsZGBm07jtvteIazXQwbq3/hKr8nJki+c3drEwq6uKLwa90JGcc1/NClv1g7pbE3zeqGEAbpA
UJu/tyBvRhYdfGFJQkdssuDhzWwOQ2K/kfKfEZm/Tv/2J+6G/GnD5KtUr+ommc8mbwXXLcCGXtJs
HMPsyoz8Wd9Zjc7Rz3DCKbkXI41wZUoP7mYgFuzSnB5dAa4Wu/f6Ul2LypGm49Rpxr/168j0YWU4
sjIQ1emOtC1KLamQ6jxAWzpE5AoZ4GSLWNJpmzlZgH4GeW/7ZhcxNQTRqW9MoRgKnb+haOPI+3G7
qxkWiLOn+ZK5e6KnytP9O0n3iXbkUwVacapgLI3NN84JNzEwvmMpGNWq/sNAWECyklfhsW/Qnwau
eX43Of5IAYmiYGbCBX9n9OR1ZArvDKJWwmSICeouLK9ED3ZhcggjMaMEOsnq3te8dADvM+Ln3D2B
n2AxI8ZfE6Nf9X2XZjLyWr5Oj57apqTx67hSmMRh9uKmm5RATovjmb3YyOTcfp9U6TDBlCZOuDye
FQGw01dCiIy6Y6qhmSSsyuqbw4n/1v/O8iLWbwCYGLAUleI65hidxlAPGVlkQuSgBM93skG0Ecz2
2Oq4uISAjcdA0wxbCppGyu3id/ATHOcYQQFs2T1Sh/2OFY5ACMKmAET0c88hbpKnkleDDj0OMu+2
YMZwY4nhzCEcDoqfrcwlJFQ2m6cXNHVHFP7/9xgYJZYqtfUtLe7TonuxOOygY2vio+oKRWopMWsc
v70Pw4C4IE0s5fVau/R7VGNESFY/E2+MSVL8m2srUnYDXFQXdGFex84S5cTy4xyOa6TmD6MTyIaM
tS/12P3mk3z2BnTpaEGiy6PZptWqS9MF0qfW1k1woK60pqz+MwrkrW5e1IJ5jfgqX8pbK6aHgZjc
MU+ixZ0mFqu6u+ciKPl9wmDsa7ZUCjEGP+3Z3JJ7UGILzz41njDPdawddljujkWB1SzOKOPF3yzf
8RTcbtFCBihueOfCNDHyUE1ZzqgrK8Pl3Pw0S9gO9DtzXY/aXd3+oKqF1wn34a2pcnZK6Bf1hPYI
ciGIlqXzVY1l6PHe2zl2X65QizIzoC1ZLI3onKFey15IjZXmMyhnpqq4afTJMtZxYsghP4vBCinZ
EEmzs8RwEwNoZCFEBOjTOnRfAnrcB0t+jqYTn17nxrGOOG9aMFqBiDwskiebVKuygnw0sPIUnSU/
9znDAzDcNT7U+mRnEqB+3LHSxsjm7oh8bAATr6bxNZTCHHKPV3JgXjxDBqczjkWCSM2C6rwXmPC0
UaaTJGEeos9HE7xjSwW0iEPECY8EJL3kmOOxR5kzLvEtACNY4eOTuYsqWR3jVAjVb/BJODzBgNbK
IjAVWRnqAaA/cePAce4D4sxQUxfNZLQRVb/QMD716GSdp8yexIP1ZBbxWeOWfk4hxkbMxqK16Hm1
1dYJSfHzA54GYnPhYTzM+m7PjU5lRJit4Th99cUj9M/TERCatKs9KGHDG9/Y4azSLYBCstC0187+
tGqaPj/CMyigZzwAleUDFXB7KmXVIzqTsAaISDgn33qOEbMkotmEUMU6Q29qHXLP79C398weyrcN
ZYEpAnSc515kkBqgiHoFqpBhmU2BAXXHbsgeHU0eOaluDTl1fc0zET8IWAyhSluMllYJuohkIUNm
dAyMrLYk2igks/bXoVMzRJlvhmz6dI7g5cJCbk+r8uZBCyYLBBeOWclj6LrMKoaahrWJUD6CJKik
f0IzeBUZwwUVz197+5L+X35pxU0vaZPudRh20gnv3AnC6hO+MePSZNdpltLxsY8azlnGykqgqZSm
EuurZJYBqJYjkaPgHGaP0bSlrLn+HA64CVYjKjnZG37vRQLo5BZ2q0Odf5bO8q5F92P1ttGHShz8
5I/IbVYziTrYpduqyO/fo4MTzrhq2DywXhJz/5CTDMYDChUzoASRjG3ryHyJf6Ajm5vC3LUbWbuw
WIElOPl/Of6+bUAL7hhIBAVEiU+DnUAAJrv44iChzsmKfYkpRfp8k/LAeLuCaVkfNTMXyjQ1Ma2H
fe2Fpxl/7q9BBSy+xL2Hx3l4CR4A4ddFT7VDq5HPN6ox9rdB2Y6r67s4q/cuSmAbhwBaIifOCsmR
erS0GsJkpuoY9B51kHk8eAOXREvThlxR8WpSVNn/FjryvA+X6Qny1sfffdQm0YWyEFeigfD3lhLF
ycd8EqUefu88bEVzR2VyFxPvuIsctvwlo9tK7t8K3qjwYXmduB5dTyWPC5fhSue9J2HV0GAPHYqz
yV8L+Cob9+I66TjK/GnQxUtR9ZihvuGC9otH/DN08spuwUpPsjtkhNQicAJkVMQ272TqhPOVXpqG
2TVuRdSmOQGJYlVBKS13o1lbTK2Np3KYT6/QF6biIr5JWyVAw3O/D2i7Xyp4zG37zzPdjMe/iYeh
fwIIiuqjMGEA/jJG1EItI6Tqqv3MHceV/4AljeDPEvh2wXHg5LSQXEszZMB2I2f5ADXFcQp/eqz+
8mAFdDtZsvQ7JM4nawJWyw59SqDtlOzNmInshB822tIR7AG5DHLNExIYVlXqnRHTczvcSiWG8kBD
V/V6B892AYxZ1CO1gqziJmCTcorr9aKJnBUsUqQTO5SwQrO/njTiCee0ns4RRbRD+vZYUJ8ERwS7
6quTob79lSo1qgCa9G3lJ/aHGYDHmsZEIOD6+9y9GWEfNW8/0Yu8AI7V2IHYu+MbxPZ6RY8oXHb3
q2YK4UxT5TghC7uYZ8/q/E2Az0s7IotkUfkzFUe06eHDz9+MvRqAfaSHP8pJIprkgrk1rmufXt2s
9I3SlxC4csD77yS5V1an+7nM9+4oCmDQX0CYYMkZuX5fGcNxtqurA2UG05/vhmQ1H1bLwOHN8Mbu
Xh4a+0EoxMDntudk2rm5oZBlTLWkgqyPmllPOal+bOXAnP9XJwChxKqil+Vi0VrbufyMW/iKG2jt
BHC+BdsNVq2V4N7QTCsgsyaRqVJi0Vktzb0qJxXtK9oVrPCE5m8bJD0n8ol8Vf3YY+UsGdeHrHpF
dVag1bNVb9UJaf18RFG2hyNEKhjQz3wrAQ9t34C0YVL1dCoZwFHe9aSAcA3TbVqPeS6b7JDbqAg+
3BLXuT03Ai03FeD3JFpC18FoDSxRRIlcyKA0ui7mKIPWwXWVJm8NidfCTjyyqMQuS3wadM9gRwQz
DJFBongLdSMQLEs2pRP35sSsdXKBgLvevEtu8jFhytlz2hQvnzvySbCuoyReDueGmL5PGo3zJ7ZI
Tx/fKX1l5jWJxm/AT0gkGz7UuMUoungMQ9ZcqTmsCAIEWmjti9Rf5LO2TCoNhVgm5UTYVmiymNOG
bjqyXAzOwOGjVDTstM+9tp496rw3wfFgEmQy4+nhDmiMFwVwRoQGhPppHCDh/nIomODn8x9Tl08E
xlRHbKrAWqSUjO2eefJs2g47qGKWl5KxVh83m59mNJi3EwwRwQR1jFgmfSnkddNfJny7xOqvhV3q
TpKjFM9Hw0+cSfqz7r0xwkgPQDWLyVSF4VCXBXJK2Ub2RwMpgHCz70mP2+CFMnTd2Iso4fmzNPYH
C9pq1okAgRRUNtXdfub0yEUS+9v0VgJpOnv+iudFyGWOgmLC8fBlHmbMQ0mgpQikerMjAXuB/OFO
aPE3UehZ5igfeSa+gP3LYAda3h/WhR7U6a2YngAJQPzNdAxfbiQbSoBryFg5p8dk7J4drRm+JyzG
T8/uyH7uqY+Zk15OAoRjqnH9ubnQKmcpX6yARvKjYZihIEjIu5QJAx5KcV9gUrkhzS15JGXLXHh4
0mAWwuj2Xo38jLFnmKa+sCsURzorqOsoEVtDWDsz7Z5l6a8gz/HhE0sXUx6pRFbW0FcIZTqeI371
k0bv1UvyKlmwSUMxb/Ynn9XRe9hfUu0Fz5wleODzWDBc8TwUdlrz2VvxHxXGB2WUxqrZm1AFu9oJ
ExmXLwSNxG2ipxV+D1glLmMwXD2ZvFw7tE7Ud8iYtQnMdZZCLZvSUnCTDNz60+NYCaKjBKRLC7HK
A/qaKGcFlCfGgNBb/mtbB+2Z0w2LpI2JVJC/JqDzIKzzhN0RkQfZvv+Bn64SFlegBpx2A3TB2NUI
enyrckB/I/cWmqE/7JAnZJlbbF8rtmojAW+/WgabipZq/tv6MiBk2Q8UzvTWqnJeqEqz93qjnnwt
dd/ypyUbZngo9VNQ6Ncs9DTokxi3QmUMtYZwMqQzkJarpPzM2nX/zGE9d3X4+JvhwuRPkMbbPbvL
7oIXo+8X9fYQIaWsGfHjyQddBEz11YZP/SFfKOpeXZUWkiHuFAqntauWevIX0ugNsIRPwUHf9DPw
NHkz2PtOxZiKYjiO45LpO5/cxvRq8TSINciJlSQ1UmP+hDRpfDc7OWkPKerCSnQcCjpipgBFOTce
aDiWa4F6oXuagpiFjKfOTor94RpejdZl44+vMBwAKJ2awfYS3ktBExko+tMOuz4nra+hG/dXDq0S
kMYUQ8PmnbBiIfZ5TI0ziGI4lZKdyqFV3eRlUTwEWOLx9l9y6AjsRL7tlYQ3EKW/Sq8rUYcuoj37
UHi6T0RiN5FugtLwe44lSMEn7D7lFQMNZBKEcng0ZHUrq4Y34TEWxW3rREbq6jgS/c1Uw61iI29p
9JUe86sVgFmV5w/RfFEG8SLffypWk8ZcsqBicdAN95maA1nAkvp8GcUE3sJEye+idij9vrBrUQ64
0Ww5LbmuQMDboQoJacQ/SRqdMOkXEJrirwkriZiKiA8kGZkF1rIWoX2uzfqXo2PNsX/74MoZ7MGO
Bn4D0zHB+AaFW91JKOgGVAJY6PHj9LUGAdO7jOGn0mO0R3Y1y3qw+50f8EHG41DlXiy7iL9RKWOA
yN6kRFPt9oLI12/bX6mwl9KO3OTW4woBh2Z5yNBFcGUn9oh7F4Rl3pRKCpX7uWJAEdBlTvlD1rrI
wXTs3bkPnQVJE5rjLK2sHsy82Z9WgPHjdyLVYLk/5iGbK7K3uf6aKmPHlOKf+JYW5hk5HDkelALy
BgZmoF/XrrljOun6sRwoKmXvdS3xk2Ft4ydrD2Y1H+e5fvwzwOy6O1uv6EcdeYtj19ectirv+JjM
3XIx/Bkhlda3UPOQRKOYic5lspxJ93YY+LmwQsppoAgCLtvRO48EdwPfwXoXSmgnuMt0UNbcYw/c
fyJ1jNx39hEvJE/fk/7ZUWqzMiDcm/VEEC27QkBGUB5eZx/mOoyAAqYM2vPtiy6xZTNYOf3xEbEa
l6enApS2maIKQF4Jmv6aO0MfFwf/iu0LpYKU4T4AGwc/Jx/0jHVJFHZgVmQtqd/ARAQgrsIt0nG9
sZn2s+sMwRoOzdisz3bi7fLzcwgNlj9xjSaPTbHhOeqHjKyK1xYBohgfYNhTarxezH2b9psEZjlo
iF1Un0JE7+hO8uKYTXmTu2XFy7jtIlw0pP/oBufoQhagWRZDSJNMD0pmB7ormOlCwEOr7qMCMzJ9
2Qz80K5vEJV1/ODbo74wZkMs2uJ8muYxefiZoNq4ZJoTTDgTCzEic4ug17y4Jj2+ZNuVeiVu5gw0
we1J7Fu2UNYCP1vr3vcDN0FlVcil2MgpZExxqSKRZbVyJgmqh6W4ufBwAa2+qlAA03SQQ6HlV6qf
MwORGrzxkp4Mu+a+QH+ZoyrfSU9D0WYCsNoPhuf2g8Ny5AmBkN3zfoZlSYL7v0PpqhUa5QBNW3Lq
UtGNZ58laZm9/esrJslUyv8m+jKWSuNYXfZk3LUd9+Nu8rJfJ/ic7YoK4/mMlIVUJy4Bt5Bill0t
cAg1BMgwrgrFIyXxYDWKO7He8r33g21E5oy1bQDNnaZu+n5REe/NuHOOzMoPNmbLZXzp5ceKx2Gv
1TJYBqbtDEKjQQdz6RQSWQulZIEWbaJZZa3+KSupMXls1POetCZ38ECIVuIiERHmjWcwEjdZ4jih
ZSGYDQNeX0dGPVPApo1wOrpAsyPLEV3yAn+/QrvGLVdA5+caAhCfsVceRi8ZbvP+7Bo2rVeXqBQ4
5oo30u8/TFVvByn60pZIBU12g6FPauRkboVvbhFaSUgQyC1cR3IDjvjrWby53lZeGlc+ZnMsx/mK
Gv61ZccfOaF1wcIYE2ATKiOT+enrb1ww8WHy3FP4gncr68xEM6VooWOnVFgKJhNFR+SoCfutmW7W
tI+pjNcV+M6nfZt145VovuZakthhwOat6e39Ui4qyB/OQrr1qwbyRHKHTiPgsojXlsvW7VgO37OC
ueiZKps2hx9agTbJIxchVXMfydI4cR+fcMVe17SgFy9iGUsUz5tesmyntAsc0Kv6FAjyGtC3q4Is
Q3f8JTmItz9nZpu44h2zvzQT5Js52DybsBdqvp+B/2zba1mH/Rd9SkLNmj06oWVAaCw/PnFnYFBv
garGyUlRkxDsI93wncwSJsaz63XbblXgm22+gA139rcxMxbHgrYZiL0/2LaNu/mtHnTlLURxjjj9
BDj350P27BiyPcYKt5Wh3d81wZpeMvuiV57ntpSPrM2grtmbnJxuipo4hUBQLpcyrxoKR2hR+4JF
1X3iMGNBR/P5iIie2rvqR/BUWLIqMlLe9GN5tlGeEUMnCYIACTmzNFA+OkPw2HF9uDkJPaHzXVj5
VjW3GZH876i/7Lh03qSBelLquKksmBVDt5UeHVBVqHVzuevzUZEivD+Yci/JxMb9IMFmyadmslX5
qutsAIrw3qaXVSUk+Xds1ddDk9ZWowqO2Jyw1eztN3xM1ymQV9U8nuHmSroc0EJLppnYbdYhWHrT
75o/CwO8OiIQ4uZwIir7K9VFdj0N/GzQrJHIepB5hIT04oBTWFtWlCVU72pLh9+twNUBYXP9VimY
Q+xyQJoJLDiTsdN+gsGyGlJbn8Re0xqrmzFZMoOgDmxPUxBuU+1BpG7sEm6dwN3oHg3HyElWUK0E
+o1jy9rtovY/4Tm1/eBImbGt9/9HFZHMEzkFoKsSqWpGCzSU/xRjqKPHdD/VKVdk7W+pSI0ra+9r
oPJ18O63rvrkjCy0OfJoAukK66uTTpITv/JYtKS8LqNFIDyrcZrUNTK+kQb3m2v8W89L+mR32ERH
CpBDCU9SWo2RuiI/oj/MSlogwPb8lku1sSrpicCcYLVwnHOu5HgoPs2JymPMtQTa+vkyhvKyh5+3
JwjWCKoUE9eyNn4n2ZRDUSTmvwFMbUMeaIwVIzqaZWtWjXgX8XF2/Z7yyFBrrPhdh9Ue6eXBLvwq
9YzDLaeZapBl5zvubP6Zaoo8CHN+3P4KGIeSQ22m8OvJzfT68ZJ0gCpCKPs6ASUalqc5wlufGVqb
mFWGTFrjxZIuuCRNitT5dmBng57TS2d/NyXkOqnB5LIJYCfM5a0zDJHZMCMlui4Kl/jo4dNPIhi6
ReFsb1gfwspZezIgA8aZUQbWgXR80IzIY0lv7dPyLYzgNGqC2Cz8MIrOn/+lFZURy1UlU5pab5CG
4cueCG6RST6MfxGfkUkxjfO/OmLIxobFP68HmuxVzVeKkZPi8HR5q/j3TWgLQKx72zWI2jplPUjv
agX0KwEP9ACsu96/6yWnG51xt2KIDO3P80DfVNAfLaUTGvxquMJ/CCT0qXhTKYROvCrOI9vQe3WZ
2/ZCN13SU7YuATL/1JXIlg6Lm/lD5tYPlQQ6ZlgSdtNxXFcI+6lQVNvpaW3rEBvv6yjvYGSXFcDJ
5FFnYWCh6VXsqNh1XJrgsAA/Dhwwr9QH40wSnAUZUp4lVwH1sVz+LK1CNa1bqFJjVvU99lgYBOfd
YAHHz21FbQAN4uQ/oVuyZlMDzqQn0lKjvqy3361SZX188ft4Pm7D+wBnGy5oWF639f3TeUX6mCMr
YioKXuEd3rSS9mTOHUjL2vEu2wcxFO4zv6PGvW6UPaQ5CZgA5eBfFe4L9BM0AvF2d7sXlyhYXSi8
brYBSVrRcZmN5yVEFAyIylcJsxhqi2rm5amaFcDztyebH23fp47Z/dHjE8z0dAkEQ9Xh+lTBKDcE
s3ee1RLGZ+LL+idcsZ6EsnE2BgANUjXSSIxWD1Kv82bAPdMPIAuN8IIB6etKBwONtPEGvqD1+pWi
slQ7aRVpCNaRK5CE38ghSW9VouEK8hxaS/uErsFG28O/lokx4FwnsxxD+apFJgob63MI0ZAX6h0a
0FMUIoSXRV4OfSLgnTZm8gArp8P4CYO1P5/eq7dXjEt+LZrIvKHbpmxVo9CkEfLFPj2bW5FGm+EX
rbBVgud6L7NQQycK8QiMw6T8nfTsl3FYpWZNjuwaKBgv3r98cdk45BgHuRHxferFueHIg91lSFTQ
d7oW1H/JyoVOxOgDSUHuzGEiOJsbEudb3xiBL0F1NosHBMkEak6Fgkk9ugq0JY3e6c3oi+YBB1du
17emdptvrNHZfWg1Z1DAzUUnGnhiTcVo18HnR837catKZA0tlVYm6HF6y6YDIj+fQUQ+l2z0ptco
LJ5i/Id45r4sV6WAr5gFb0GzmO2Wi0Wsqlg63Gl82JmopjQ2KbvBN9kFLOspr4Wg0wemKvv34uXg
BTFkkHXgT4SXubMb0mVPPAdI2N5V6QW7jc6yH9d/Zms5ADljPo5ocoyCQqFDa4bUpc+yj7qKdyW8
0K2D7iiNc08UEpKluWFFNB8jAoi28wsJcUIJUraiH9JYvu/k1x8U2EP2kLKcri/JFyoFJ/Uo9VJg
aDAuRqncO+TsnhVHn+lAWHj009g+JyjLEFbHAcdHHAtUTTOL0Li6TjZenktHZwzGFD/6ztaeaAhA
SSb9QCKNQHcw6cvLXUzcqzg13CtcJJJv33EKlKEYc9xf0LQV4V8BvMtm2jpt9eO6u/Cr2+1lg0PF
Nnq7IZLpU/67UKd14+IUFTCsyW7I3On0AlNSrQOEoVShAfxRZrPC8zcQ0TGlPxinxnINCKM9peTI
uZKzbesI0+J4KOBKmm34GyjLtbES3Chq+icVd/LCdShiPZg50Vgp7lS/d14OccxB6rp/l1EU/zZ5
rcjhSP6ZqvXB3flzaAuRpZZBjZcS5qD4urIigDP2aE3psTSS91WvfnO/OHKOcBgx6+z/YUMRktnO
G1sy6OfE3CMTeKcU0pn8Sda/tUCkQX8AgQYrUhWlrTNO3QHTWdDtKxbv3YtsQGirWcYGFUTXDpiL
WJR4uRFLMLlEd+znIsOjko1D9bEhsJUXGh5vKfuy+nvtbFIr810hwprGh5clRUmqL6gOWHDSXX75
XTGsywEUV2vYMju5qW7OnBc5XGFA6G8y5zz0C/Tbdv9XJDq113AW7XbXTMVOviRSparEmjUrlD9p
higsqzv6k5pyoLdv1nur21BqlDdFTSKjNH6F/XBB6T676GlM9d0bOlQ+hPAnmejmBNWbt0gct7cu
LP4cPFk39UkUp7JI4JzmVyC92RImeh/wf9pAQ2CMg0NHnnyD/J1AGjaOBW5GeQPibxoyt6x2s0Ua
grydTc6J33gvitMzmgDDfTtCFexTLWwe18zm1tK8riDf2EVeD+q0dvRh6M3INqVGj3ZSFJNzmVcX
xSBQCDaQH2+SWQ03giN+3C7NV21/1g4B9PxYM7h/AEXjgguGoyeKi76F9GN8YoXoPJ/TR0ZVovxD
YZ9e7RIA7LZmasGO8VCMLGOBT8uqOpfLmky342BLZSVrLfrOvbodsxP4A8rWeOsb5WWTvCjU+5bF
YSLMGNIJli5C71ZwfwMmV491QkFbG1Zj6Ty13oFOjwYrIUl8irbwIUG1JcMNgEe6886JYtRo43ud
REHAqf87+xz61/o8XH5mhBCaSlOG2AlYZK/IcR98Z/gC5f9PMFTSyWxs2rF+E0BH9FEUEHjAhKHP
DK8cQZ18a18lqJgN/lrVeF4VxYz7SfA7UWdUeeJghv67eNXLaPWsPNSXWMWsrC/A++3vNM2qE/D+
UHJnfVWFbRPim/NalBjZII+Mg31NABfwIuZDR59I1GFHNU8ZrMfN8I7NvBtQen6PlJNmxuFEPyVe
CzsVr7+7QD2dYcK/KILkQoqhCfT/tQEch0kFDxf9am+VL53V0JMTAutjH7f3r3P6lABWwDCqQKJG
y9CYYlTYorM5ysj3Buwu9Cn47JKq7aUXu4U1LqrDpJ+UdWIfJ5/FOpepiaVPHUi9fWrceGPJpvIE
uOdh/wxyA/plQikjBpKy+6hU6dguXirR+I5DJDVfyEX0r6klfKmLafkJkExxcr2EXn/UmqSmwb+9
0bHYVXGtmKJUoxGJYZkqF64dl5B0IAvyiTkECuUqwDMfpnO7+Se7ET/mmhX321BTRArdvljQ9xaf
oqowH5H4LIETrfD0B/MoDKmv5GXZP2zLjAon7ScX9oGc8cUqDlU8mtzjtTkgBc1+SKpLTkcYYBWh
41BpS8/UYKYaPb0KeXNuF/LHsWTdHLPIJ+IPhO6yExpH1z8WJ0+2Yd42AvqLCtIp7pWfJcL524Gh
iuhhnFU76phJiYDJf5/RmlUH4K6IeBXFb7b/t0My1oXp4XivJT7z72mmELgIiVPaPpOciG9f6ByX
tU696SC+q9PptlC61DNjI79XI7fWECFML2ansG30tXY+tqlZKLY9LIqdvSsFIN/trsYil/Akq5bH
Kxq3qIbrJj29FqfcqBXmQVPx3Zn3Zhsnr6pAsBp9zqHHAQaxLrmvZRcchL87yeWq9r1tp/BdGQB0
heXiFaTYvfKaLKjgvb3k0Jm1Ztzjgmk8c2mN6Ci4HIFtXUKQ59VuZbYRUdTAyHj4myyITUvVpcpS
iY2pmQUJPXh/kROhfGnGv48KkEkD8lWrJHSjRxNEzuTGK5pbf8SOvKzNqHKSQeNGsNL9ntFpS75Z
axHVhfTu4OUFgMMx8AkaYKYB15ac0eX3TQaZjDSzWx32oavWy5zqD2M+UX3vV2HbqzQe7JQnixCo
7hiBZbN07CcSdwgOGFC4+/MnGeDaDk+teamEWEGMtwayzhNSi+0roi+c8UpdmSKbsNAAATBR8eZU
NhYhznr5+7yqyUd7SfL79pxU+m4JdOkz+XO/4GQqX/NFGGLg+U1jz24Vhxi6LOV3ZCTCaD2QHVgi
0S0otaI1CxiTnR7spg1ulDXxBiPyVbGDr/vgYI+khcEKk7q6VfzMpKUyNiFnN55GDO6w+6Hz7l85
Wo7b24CuWW+uwHZqL2VaOq5wm+VaHNUkylYkk9hkUoEd8LHIWv3IgbRk8A8bmFnCl89Z1sCwGIJ5
hCe8xK47hlPMdfN9KYqDwViFBUR0cLJLNSeCIMeBVvsdTPXZBkItfMDcZQvE0J2Y6ynz1jsOSJ04
qpw2kHu76ZtG8sffNeAGW7Gy2CuqdHIJYtaqz7+Db+1QR1LCL6fr9QYUWTtt7XYgmKnr0n8FFAH1
rHVHOvd53PnhDPozRdxAigPnh84Atbf+s2KKTaHKN06rVvJFSB6Sm5Eo83VZ5HLuwQSuyQrtIWZR
BtrDuFoh2lvlcYh7HEjr5SzTHBCLk74YiLdp4hiCxUPpSrYc5BJx2xfwUp9Q4/7y0non9GwAy0tY
Nn7edJMQZNPQU6q+I913w5y6UA1QQNZD3yeOaaX2G9d9ZH+vGej+0YOUdSVUMW+UVkf4fJLqGcsf
nbAPYn5u0QbsEMV29ILeNlHvRJps7qa5MVtsR+6FJxL1v1F/Ev3ZbhEXh37KWVXTisJbuC2EOkCk
MOx+5YUupsveanSXWajAQhlc8tbQpVQAaRUjs6g12hFeeiixFsI0zY31bvJz0jqk2eSOCj5tfnJl
b/KJHNjk5bAebanFUDQVM3cFTiK4j8XHwzja3TTZ0RRItlWgwFebtPu74U1Wk8h74UmRdKUobEYP
4optxMOEmsz1Zbf60oKIT5cykOKKpEVi7NIqzo/bEoRvsd5VgCpGV7poTrMsiGuF4u11SaPiPMOV
f8zP0v0JNxmH5eST40TIRnGK/RMRpCqhKmVZQ2WYrhDKs2oom9W4bvwFvaPcjnFL7LpKKTvTOpaa
JmWPDlIqyhfqKkN+lt+TRYOYAjmS5Ai2zy8pD6BU1ffvae5coZBW0bvz3WnyOglkx95tyRsUK+dc
lFiTwi/M+1zCE4K/zvjrJz9QUDoqgqjIhYQbVlbVTw0+oh63xcofoCPc968ahzq0Wev7mS/A+OBF
f/ucYcr0uLtRpejpdNnJHIsg6sOT1DHiDGoFi85Bqsjloy+ql2EPLuFqzNt1wIKg3wXuKZjwfYFu
mwfWxU+vQczPNUwXcU/KLCqXNKTWx0I8i31IYimk4vWpXssJee9CKGVkW1uz6/xUZjQLMZunBsES
qGSZD8DhRWgCBPMZLIHy75VBxEuaskgtFuJSeFLcGHm6VUYQnLqk8Ps6p1UB6txI3D9bMPvSkXE9
s8kUvvsURg6maLOzgIhvBencZ6ky7gLXSVKlkA4qx2dTg7sfW5ZBL1eiEFTHYZpP7A6JjDKbk9//
WR0ON9/E3zcddduJ4CpvVpZC7Gb4ICnoKHefv2+flSzstipace8IsMA59lHidW7kgPDhIEf7i0rs
EID7/JfH0GljFvbH4IY9yJbBgtC5X6BeHAnAKgzCKIlm7tONMlmc8TWHwAcRYdM8WcbBwp3VWsVA
X1k9wqZEdcbW7Xjo7sdrbUDBkp2XgDH/h1/yyqSkHnvGsUZZdyOWS0vbzhWi6sXpWiPCKr+SNRQ7
OrO8+Zwh+sL4VFX2Za2HcFs8fMLQbtIjewYTPyjFOjekYcrMEz1WFcZjnK6UvpmZAQhMV+r+JtYX
QUdkUefYf2IqWRQmDiO2EPbBkQOCLmFP590MPV99GGogSLX5hTCFAb1a85mDnQ2HE6khWpibTTEY
H1cC0qRzmNjY7X0UG9NLe36nNVmdaiICjJOLE9HjbnDd52Vfz5iTZOWtTJ71tJmI7cBWeIbT0H4H
wFB8uAeywaTSMNM+pzpCRDvhBAI8wPpcqjE3NbdbUtE/8ie7NEmpLy6x48RhRD4JVnShHafl2TMA
x0QklT1U5WyIGG7EqowWB9cCczqLbYUa6sWA05Th3ckg9ZgnR4/g0KKmVwcvPZLMpL5RKZryc3Pq
sYysZAhBcjY2anX4p6AqP9J4VKBoU7sadnxNTQ9we8SjbvL99TSVkbqUgxzMNcEJ3RwcmNuReSb4
xtxzrlK9ea1kEa7xn5NXiqgvfjMCtAkmH5atKAYO/Si+MscY4e7fUCOwcxj7kTseGGJ4upz9a2Nr
yLfit/zKltAKdsbzp3iIhz9O9FxYl4SQM/M+HiFYlxopBlT2diQ6+vv0pgiKr2m/aX5q8ZQwv2cl
M3VwB9KKS8VYmP8CFVI/rIljg3Kukb+M5UTUALU/ZlSd1uMDeARA2sMyETl4iGhcJF6mwywGA7+S
08h5Sd5QR4ncEw9Q2UWniaVkhm6LWDvYGa8HBY7q6QwBkzjQXKLRzFBIr9dW2MEWiiAaWeipNi5z
iQojadmCCEklWokAayOZLteWwrEXnHdqharWqf0WSkO0XPPDXAlqdUG50vZ6DafWqAdRnmlOkrnB
6xsGlcFq+/48q/Y5sK1d9Hob22sOyHK7cMjXtzeo3kXNCNTu5rNibCgswAnAJo6APWeWpnKWeKKR
rYEzD+e2N3s6PhwSbE/b6hcdvZtxDBq8+CRphRbxpAcO0Dmiu0OEoNJSCrS5FILYqxaj7NbshSNG
QiVrPaimdeDZVLP8LlcYNyeCnEO/5X9VYVePWq+sdlK5Lb/maszFk81PVVLVQePGEXOAn3iA31Jp
KLY7o+m17/HFGNRHzXt+d/mh58OXeSXnoK0+qA3gN7YdwRVFri9cJZM+vgbwFM+34p+MVJYjHolV
4SC4Tixl4ATyR3QLgtFRpkc0LV0JDA609c9y70sYNKJ3FkEGkihSQrCb7B8EwB5xlYkRdzC+Soy6
2qlnyhzyT0yygA+RolPGFQLYoljmQMq2lPqRWfiO+QjBZwHPDLsPU9CCNs4EaD2ujWUa2gPEc+MD
iWJ4rJpU1o/qd7jw8q65UpBL6cKl6c9Uls7AIGmiT/BrK8VM3BDsXnS4dkrYAQK1UikzAqTsG4wL
XEQSnjP3O3mmgtrCGAcupth+lOiyt/9LbHe2v3mlu6KuhruLZhvMsNxWXW6SOM0s01fUYIbD1UBv
cmYADuLICg8T5wxL4Rgpt7oenoU7QOdkzHVHjjvOQ0gPFjLKKAmtBvBvywothvPgpaYb+PrmCxc2
0AMhMRjLNzbhrYJpb55DQSKvSIB/TwZsy+cPRva9XtjMWg6oXpopO/rAVb2lrDlP8aENgotynZSI
vbvWE+7sYJ9YlqN9VwaB+60pQm1GKfsa5T7nlJg0p6IUlSp1R+YtO2PNrUa6GDn4apRWBorcCYB1
2tHRkdpK3q9cq1Qp6aMPRxgYeH4Kn+eougATbIh47gjGYtKf0W5nwYdDXTmrbCtFXFPnNTX6Uz+1
E6bnd4zjwYY9/Yik622teDSp0H88eVLurgwIyOgooEtO7N/HV3yEd0BfIOPwq0nbeqIIJCNxaycU
snUuI6oUFRiCx3gm5DVsxScrTn0bsmbHLxU/9ciRigUqihlMURj109Efg53d4/47RcEVJZHI1p61
1OxGV5iDYL7nDEq7VwmiOh0TdZPPzcUY1W0wpEuIp8Px6CKzJviyKm4Vq8LWokfqIFxVY5H3e2B1
94daJxTOQOPQmzcVWtVgpwPdtsi6kGNXxBh3qt+67Q4RtuKLheQzU/L87GHyh3psmxaqYmg56RJM
jmKG9JE/usgrhW5qox2RdMdirmyVCzQKoCrVGrXYBNpr/jLRw47L7orpFg2yoGZH+EHQU1/CjfOQ
99+N7xXcIH1f3yYrNbqGkihWt/Vu3TGD0cvOFEgK93SanoEXYMYUQg+9gaoPoBYJY9OcYdNc10bP
MQBygOo8UqIjq5Vy8ObnrEyhybV+dld7iryCn5YCkdUZzXG4f7WiG4eNgHkLmXg8kHdd53gkh5pv
GOQ1GmCp85sQPyDALI1aqHvYmIl20iHPzJDhxGWi2kbgG4hFBgoOqhVBbYaAYbRW1VxYpgQLbblR
6Dt5SbjInoCmiQdYAN4lQYSL8TcLd/Lzl8HBa/V00raZxzZvHuE0i/xWpNYmwuW46V36375dAehO
gJwRozib+zmtX35rWRLPdHg+ZGGzvLyc6cIdZOeLvIGHTBUh6m4IPXhb0bD8sqvYgbtHB8V7qxXY
HdQ9cTNYHZ5e5Snwzk+dibj6QAtnWWzuRrtbvrIQssQDqFiPZxlVjBoOvsi2fB0vkrE80azoZ8iL
BhK+S6t/DUPfNPwJcXLckGfUJ/wlPuEwQ/XIW7Wj/iT8yURgmZWWBQvyx/vFPU6xeTswLFGPkrcC
hftUMGcNpKsCsMrmfj14ErQ85ybTy2J3VrQ+YHF6Q5PNHXymaNdEQid1ZTBuPwshEfsa41UzSwKZ
UnHGYrsFKoqevN4yJeSpEBqdAdPoKesDs2USqjWvLIOEO2zoPRKwOnBV4xqDRpyhozbRqZwuNPb1
NMWjK/5v+/bpjeCci9kylKkKKTq1tKVxGWu9kxqJVNZIvc5jEr9m/tWAY/FGzRx7lyGPJnj4Kldv
0E68PEsGwgI6/ni6bNdT3M79xVOCSF3DeuxZGpJ+1ZMzuyxw13XWHGk19EfUg1pdk66sTXM2GI8H
jxJ6dtEyxN4FofVoX+i1wTebJgwbgzN2E6PYSzLHrBaYMowuDSDl/Tg4KiCazFYzx8BnNmSjbg6F
KgJFjPY4HLdY9iKXTdKHkB6AUG+FxOUTBWt/DJ0Wl2yDcMpyEEI89+PjVfoeEAyieJPOewBl1/Xh
NZijs5ycRlnUo3OELGLL2BuzB9oKsjjTLcOwENvUnLPRCZFb9J2p+N+gUanP6wj4vBm5YT8uIxRE
yavbUq+eLIaEjyJQ2NOHB0tObUt86a/7ILyPrNw7Gu3p1XDZmMOqP0pIG7JA4x2zy2PS1LX5nyN1
znkxic/b1iSHVNMfSpmtrOoKvL4V+v3L0hUN0R3yjh9LdcnVmiYBh27AhtCWJ2mY1f4OaVf39Qh5
R5GQE9Wt3sEteIDMahyBD0OlYQttfjxL/pacLu+0syjTRTPZTP8tN6BeH7qrLm+C06A3Ac6fHVcT
ne/TVqvnFf6QCcpZK03yDyo5dPtsg0eSfWJKm60ZqiSsKey8bepD9bEV2eyEiIxHXb/acETB5sJI
FDFFsWAFwNR8gbbMhiV1HAVhtIpzrvpv96euN6/t7Gs5e1ilhPIn+otYwVzzfRXzmzseyXmi4sIN
11HxurJ3iVlu2NuM9zwbbHbWkH/B5WGZLqbSuFEbP2DV3R61vUhQRtVIwBnxm6JBh28UMjIOAYXM
2UYR6vZkjg6eXrTjGp87RJoxXmkGLyTVzMMsVhwNt7QZDBqfWN4OmBWgt+SB/u0VUfpuiBgNBsDm
w/fxhOYMK9dvZqECbxJr4d5La5/Rrm381UoLV/viVOqXf6SpYMiglgUVQ7BpGOInsMFQ7L3xPsP6
y3Z0EObqN3i4K+dVf7GxFcuStIWts3Nvtf9zbvN5ZBI6L5QBvGOqmfy2VdE2DnMIZBKDIm+wMM1m
bDiZtsrMYpSVq2S3BsaNP6PD8DzasdRl/SyzaaqIzsURKe9tjuWT8HgRj2MowoSksBqqfOA3Av2Y
95LWYDumVKuqPueg1quFFmwSTDUFmv1CBwhzjRRvBWBFtwg9qzu+hToBff+C8kaH1r12kAPujf8s
7tr5nT9qcmTUjVO3AY7YHjLl7sHOrKPjG5fji5zQW9QGTLG9nNGShM5BsZH6+f909GXxPNtVkY7h
zOv6AygjtlficEbZ4a+8ny2yDzmQQL6vrGiUcK43XspvLs67ioc+mFp3w5vHS7DNWzSrs5uk8CQs
o3twHr4Nxp3Vx9PJYnqVGG9bV5fmRs4LBdJhoPK7+HsDGTmNtf4t/q7kIN2EgKLR9Xkg1dkT0uLL
KbdMEVFVLmr3Y/VxxnoXBJSDIBwBHDAatmrxVmtbZKF0eFH74s+RzmK9vytgwTaafYdaznULIjeG
ZhV/GXlKSWaNp/WtX3TvzOo5tTsGOPwskRj7HcXh1dRSnLFtDD+0Mzj14w4mkLqga68aw9ynm+IL
RQ3h98PVLl9AeSM/3wVe0ULW6vyXyt08f9BM+AShhVvWSU0KBf3DpLeQbZ/+vBZvQ+EfRsalc9uQ
Mj+tZ6BPThBiWxjq9+JiS9bb2xtmIWMnPjYGdnYFWOCmfSFgrPQb+UZnvIQFYSvcEwT+cBg0CS3B
Jx0ajtRci+sc4MKcjXzAXTZ7xxil6HcL/MdYCZ6/caZs/rnXMZjsTjHFSdbbA+RMM7vwEbq4Fiug
meNm6FT0VXP+fdOQiCRtMMB7QUTQiRSMlDE671je8zXyi6uHl3CrR/f2SfLIqw7pnD+UDSIECHcd
0lIRHRto0wZM09EHnIaPdWEWNgYJeJwQGEvWlg2dVGK6vMnprAftrgcZs3t0rnCq5Vqx4W7oKaiZ
7ATP7NAh/JY/3jBkwMmN7sbhrrQ6fASyxJYTST96kt7bZPUVKEICVitar0FGP3t509xuKZ2GVYlk
dptvxtCSMg2q1PhlxeTgxHYeIK1nTn41Uj3Rydv+EKzNAazJmiJmuR+o8j7L9dYszR/KBOJogTVK
8I0HDIeeiGZ3tttf/1OFFvV3FG8H4cAeh3bfKttGaAzr15G2vgWsB7Gjmp4Jgz6uJj8n4GyfuIZ5
xNmqje0rwFN4HtkCbNhHlmzLrZR4sv1apYThpuJSVf2LGbk8zNAntTofYitkPMhsIMulmwPg/F7D
klcg51rwI4EvCBfH+hi6Q84t4d3egOya1fkLxXUlubOybsRKpeD09dK/XjBQsj/V/1KStM2nzBsK
czs+LM8l790Tnd1Ln7s9OhfT/khdjIaTIxLh/fxTodzLLcYJj0N1k9ie3gdDiyWYEBphBWwO9xNs
1aqX3RJhxGZ132v8jc9cYoSdoAqYCEDhjOxSl2RaOzO+MkcPrnC+HfMglVNKuO/dflR1ZIudJ7z9
++Jg+uDqAAzW1SyGl7T0TAJwwJhVMj4D1flaV5iPEJ2EzdnJzSeb5JaPngCMsbxj9HXZ0CunrmaC
/fKXq3l1ii/YJPT7lyu87QkiaWiv6uT4CZ0m9Xm48TbVuuPrAlwy8ofNh+SsNB7NWB7Cj2cc3d5/
qOG3oveV98tBtt866Cc+DbbDnfCuQ0DnSHcTN2B5wBKddwistVRy5yg1FKFRc0HdOr5ciSAwCu8X
6KZWHZKtsOT8WYdI5MUazdc7MfnH+iHvpPJBHphTD8ZZp5ffEhx2H1LrwpFV4DeCKMZfm1SZV4sr
o9K5W45MSf6QYBwGhtRlkwiIpIcMD9hjqH6fYFfb2LnaF6ZekWpT6yq0Nv6I8NimqGro3pR6TLio
7j0WLaqNVUEbIqHlMlAFYNwoeOH+GGckc6sVu5FTCOwiPkFW1m0KzQHqFQMhLKHZeVUEmSWdeCxw
TOJNhnCzhYrY1RfFY7QahGCiWsaGRRolNslgDBMH7OMxpNxpkGkiOOna4aplnKIE0eCZR6irfBGP
1wtrO5bFHF+v1PWn4oKSNTdp0z1W4WR/W/zmk20iOl0YMXiyEv8M5FE9QnRv8dorwkIxZFOW8YrK
HXLx1WgCihy8vjKavUNdGpNTe0THKOEjOfxHV7r8HJP2XcW4+gPN8dKx5LMo3eD41COru+lQpzuO
AwGsPPWLOyyHQpa87Uw9wcMBw8jFBZbJF9H8CACzVEBbZuyBAPjgY4Vgm63+9S+8FIbpMhsOclmx
cQ1cV5FeR0rEfF3H8WSuLeNjxFfOBpuihkXMJyCG5+pVWbM8MZzQMfhoFng2q1RnQbnQiP8XbMDU
MSDpOiTZw6aUZuLIoB0kqPD4o+0BL3+YSF4LLfgg4yES+xpDi2vI+FvJ8ZGbYl3/DH01IquvVlwU
FG43g3490Qoj/xvVTWVAw9B/0kFj/H0+1mFOx479LBNkGyS/RNpVMBr0e1LMtMV94oZHfqSea0Aw
gCe8WcZMwkfvWbLP8Nm9lfd+0znLsVg+8KSr70wD5TnSMSlmxTg/D8swDYS3PUAegF11eZbsPiUd
F3hL19bvJpNqq+0jNit++ZEscxlG9sxbboWSKaZb8GT9UYUt3VLVxbWDFAuxpN4/54Fw2zUVRXL5
TDm7mSto46nP9n7XqETG/kWOLsBTU12xEpT4YVDrnkJfAQLL7YotMN9JmI9I822+KneZrgmy7b7z
XPddosAF3mfJxBIUeKttwPOQCRlodtYhwyahEfRymAUCj9ZMUR58W6JBoBDL5Ce49yKFSIRzf5/s
AFStPEFlVeaegRdTUGZQeP6RNsPi4Gy6eL546WrxP9eQgIug6Et0Hk4PrbtH3QL96GG+BImuNfEd
UK6oLr2kK06XMUnvvG53KtRPrFHVDAmLp9Cm0/avFufMYu9ifsUKc25m2VyfgEUaRYzMkeEIZOnG
I3KLUQw7cGLJom3muT6y7JkrLFbqnQV8r+UEB13XPTjGMeeXimQLtb99G6NLgcCgWCw0Zok+h75n
cYpvzpvFRNZdU0qCi1OCNz4ns0gAITTeToTAtMsMjw1fUONTqlsc4vcGRrx0cXWwh47Fd0ErcB3A
c+0r6wR+GgMaVmQpks66InAnd8moJUmbH7MhqAJ4hDNLJHjgnLZ2jZFwSGJTlnQe7gXFzYaHnWcq
oQDUH9Se52xLrFCmNeoX5GMkHOCHcVaZXprY071/VjRoEGq/nZXJnwLnvm/t9rCo5AUBpsZwmtn3
MTDNROcE8e1I1pZjWs1uRpm7AYTBuYAoDcQgwE55jFqDxxAc6zzFtGL6QCmbu6D95kl9GmM3saEg
ZXmB9RDROdIrN3OD87hYdaeNOIHHX9eFQY0LlXKJ348jbCvjDQ0eb5LNvc1QYmBa0TVoI4c046d/
WFtYSHGg9eUaMQRgz9Hhc0q3cpXaSx7oohfMo89u3aR9JBWum9BZjBL07ufyQts67F00dWlYwi4V
zD70ojjpgMZuR7K7ZNjpwZ0t8tetG4uEV0KtsG51m6XhuBjI+dvDC6hxU0aOX80RrBhya1Rlq0O1
aO4fSJ6IBYNE+rhKfmjcZoeeMHTxDCOP+w0gqDI37Y3thmM4qeGfbJkoEazJO0JyzIlfc6Bcsa7z
EdINRkB3H4r3IVKbD8uWJJRk86IJ52K2Fyr7QZ5Tuhc6/8fO1CXXcVh6RcUB6QysmTwlN2Cr4YzC
/U4nxXM4TM9c6vKF0JU7GFoh7yTqziLCx5FKy7gZ2cT8Q36Lq1m2aYqKQ3gSB6UTFG+aSED0jnkg
cjziRhPAPk/dba7eUCvvFxswCbFpKKCbW16pcm2jx/0CHNoGU+lYyiLKVhpg2LTjnDpRf+8SQrL9
+0Q0l7v6CS03AJqwFX3uHakysZsd7OIGN5GlF599zX+gwccEYFjzlZj5SV3yG7VR3mdGGyjVIp/W
cVRcvMaQ4cLXz60cFi3vRU0p0VHQt0yNdUGWV+faBZIsimvUHHqv7LcirYudqNUN1BwjpxKhDDQf
DYIuFmARl1VfS+oDUBuN88HYYIYdbShuCQL04IVwck05WcK8Z++zjF8gUY5BFj0t+Yjc76reeuvV
h7rb8dlUYhj5cqRLJIQNXpa2ucxCvIokOYRTJCVKKHmgYS7XGv+qEM+t5RZE8GP23xVYRC+U+GfX
eEqHGwMGnbXUXGBrftGJyoW4lNXOl/uefyf9CPxt49dqSRSUfQ/dhl3BAcKgUG/WqPHR0fTtVRdI
kxjKKax8wxKcwgQD0YjYslENhxqWJ5oW3V/kGizFMdf7vWZvZytQIlwsj5SYta33r+p1wEbURvrA
yqbOfWdxE0KcyconMbda37e1T4sQDRYrwKqlr8/k08LBybea96Z6KhpAPMTMwOkivnrGpMI5xwfg
9iqJGT0jNFz4eQO17le/1K6qZeHhOHHg+2oBSN1EdshgXVz5UqCEEVnMs6F1AY/YRuS3q+hrXyel
rRQcrw8GXeswOcbVZhEuMD4Z2m9abba5qiPjeESqPqic15b0kwM5Ge50VAttiFTpxjkLCjfOIzAn
MWZkC2b6e0wRR6depSznwS0zz8eRPhyzJXYv6ARxyQuwlu6GJtSTXuTuPswR9IAlPcp7euiQKOap
zZ4xsOUh0h30nvYM/R4MJKfB203mAXu0vYl35Zbl8F3TuSINARxaWbp1gevoWKeY7JYRCicdniWC
t6k+m4tTJ6sBa6ftjs6TN4aTIfZCuy9bpyBqMdE0VwzxpF7wzPmRXobrLpEWPdwOh4kpn9twonJi
tNKyvjPXBoGo7EJJDbxAWEWF8ZgHllnUr1ESqHgxXgSHJfkTpYBiy9GFcdF0Y4luaPVM4XLr08iX
GdTDWxIrhpagrGgSRhOsaE7TRedQvEaXWwOIAkdmmP/CGzX98IQGLMa/9MT9cQeS+JSdmcPU+nl8
kJYIaxuSnqaUX/+pW1Hgw76L9qvzUkkG2LQMvmYF2ptH2PKk3KcJlglWYhclEGC4n7gqYV9p729U
nuelbEFNcVS/b4uvkejWf70EyeguxJZ/6lsyOFoyXqsKfOlEE+KPXf/6u0mGTuoM1TenmbIx/fLA
ALE3JBU2VmUKveF7fiyzcnKjDWs2Pe0c9LDu7Af0Kx9P/YeijFaE9Gnx++a2Bywn6356jDwLqdzP
Ri3iNznG45CszKYRD3kMKcjeP2bwG8py/pXRS60R/0IEYg3LfB5cPwIW0ptKW+jzPJTO3O3GAfOF
ZUZf4ioiG0uefpiGgcqtcfE2n984wMlGz6RbXj7rppV4qw0s3c24HCbdUreiPLwGlZJUH+hYJPYq
sZRWp5Ym8JclECSzS0I6UfXOKVJwHrwNyVA38O52TCvk3tzTMG0VKA/CRocysOWkjJkLfDHoOFuc
/ymYKWyOrdmILTQsTGcGscbf3NCoAc3bCa8D8G/HCfFFGHczFNyyV1GCc4KpKkOGbH7TBvqgHNJZ
P36AKuZ1hU63c9FRXMC6dPIP/9gg8EuyecpUCzMAsjVGNV2A7lYPq5Pi2mID0AtpGi9N8LhakUhi
FWjPjly/qVe45gpWzKAowwWDVIy8VlWFqPzJJMGL/FNFpr/5F0b5fWdypSgnPegdBnmzmWW2GLrw
PzjtMh/EDg4yq2f8XC3jCNLfPhZusAFu8pGT/8HQ+gsyyRW+2+IKfbqkmVOT0D9Z5SsH7sW5HtmU
dORWvXRCHFfP2g9eBGKiEI/Yo44xdoRYiLmNg5N2MlytKVAAiN4tZkaCEW2lPvykTESrquuUC6UR
RiNF7W8z3V+HKu2HMvAxP2O8r56CofIFPzJQOa9iYTMivjGgbIDcotNVuFkXowtvRtzsJAqFC43D
rLpytD9MbnMv62rPxuUKRG8KKnF1cNoFn7hh6zJPF2GVT+rnfIB73Mg16EFy6AwbYi0fTFjN6kmR
z0dgLHtIh3LWb6RpGHvX3C2tYEmyrNspg2a03EfgrOH/qUS9BYNJfSMhn7ULqphyzByn/+21gllX
yBZVJuKgocM9QBKLLiKl2JbdgIMIXqfbJ3hRiCN3sO0wbwUmuaexUip9ZxbKDPqhZ30W+k8lkAG1
uKpeRf7kQ5fjpk8WKxoKRKwsrhp5EBIUWlsdjBQxqLqYtc9wXw4yaL1ctn+by4SHjFLbOux5dam3
NkouSWxt9G0AmX0UQcBmqDSdIWjZptSQyddjdfC1mmPaRx83jADx57nOyg1hQkWaDuS2IPzJrrFQ
/ZOseVvhZUYyjh8/ZgJwf2tjN1gD9h3i9uWaE+9m6fJq8T5cnHEhQQ7VVxuFT0WEG01lGRa3aaBI
76P9QS9xUZQWhI/ctpkM41Tx6gUx89kJtec/3BSPGoyDLl7Fs7DYP9HYX1ZKqqR/V8dQ+lb8bcHi
kfFR+Sg5n83ODYbv5tKDX0EFkEBc9TwsPHgi5XeFaBZqIJZ+PBIXPuH6U0DahhbZJm38esrbZPA5
FwmnIO7ZC4FRXNVS+FGDvwA6D6741HbeRsAb4rES4UHLtqjB2Xudx7CiBOatZV717UkHZ4ZBA5Ho
VRi7eZKM4tOB3VcS59DCic27ApIw/aZPg9iTcN5V6uj+2T48al8JEQsJlK/RCBAixdHl4FPqCVU1
GaUq2DB3sw7wCLqIdujSIwvCSj6h8hjRWNWCe+66lQVteg/NgzAQaf48nbRZkOvy0xCdCGGEIYUa
2HwnMsljgj3OAr3soFIKYU0Tmd7sBerzUx7XgbQMIOLYk6CZ66YwquwqGdR5a01j6Qv13MWAawqt
FNeTvRnpRv+FphUiwS1rxB9KXj0sbMHuXPUAcz0jbe42x7CviwZW101ElUwxRI5aG9+fYDB/az3P
hx4pyMgdWCHHtOHk2yypKBuED+oxb9x0Nr1+pP957419f0UTQSwsIIHjpEVXFU+hnbzbrdT4Qlo3
M/sr4uw6AE5mCfA1dJgU9688VF/JLPyjd3p0s/pXepOMfszlwDXWx9QBsJyG6k0XM3X/vSQkEo0i
iW5BUoeNk7e8d1cbEexNiu0l7miHZ/HUzwJaIIrfgRWIdD+fpMv7VNUf52+uXzhGKaL/osvVvnts
0qYITaJN2/2aQK4XE7ULXAmJPg9jQbyKfOSGNn1REvrnYaTw/kJqh/OF/2BsZiGGbSRQeJSpmSPh
dK4nRvtaxr3uHgx9oRCZDB3WAB9z+zgvBuPBnTsR6rHELbItT1LQRnRXD1KPX3pf26qehRB/A0CG
oJZLdJQ2jF/DpkRosuoGCPMFsI26tOxNo7ObFuuckX3E8v/rLQjXvAj0yswmtTjrUwfKjpNeGwlw
/unRJTTJPmOJFZRcwnRzZ8COLD/IMmXj06GxYfPcdNCGWuSj6miO/irGn9rLS2ObQaU5taV42vCP
oEEDxSBk5a4Kby+XV89Ns7rx+9r4itRqVDksHfzlYqPCNOEhaoetANKzd5rTZkkfs3geXtz0qc6v
7Tx7hcUgeBJO8chdIfp/VMzWersBsAkXOvyD1DSlSQkpBX4l2ZuKguQ94wyqw4JlrPxe3T62+4BR
wk6I8Y2A5FPlUWfz+YaN3oy8SBcUHSeHgUTk8Q6/O01us5LUaF2+BN+TzG6S94yzY4jNEwSUvg40
rlvwUVLZq7ZMipfzsKodasCCgIaIanJeYGyUrhHrWhXZLIu5wvsK1cKkMO6++QZXEeQfzQtI8AO8
LCseQmXM3H1x2w/ML44w7276qjmqsufNV4if1VCqySmkZubb6W0U/3mpugTK/pwp+c9+h0ZDXw2q
Uq+QOtnVBkDd7mvpQxG4wjcSDhRLaCJIqzLOQolqukC4MRSs9qgXxEH8zOeGt/bGY96bBM06knLb
hkgbd8w5vmDSYX7Zxu9R7oDEv2hg/T0gnRTGkO6hEbKBVlGEs3gRlwt+2DSaq+893OAXyEheczNZ
hBKdPKQiNvhR2hG4NKh/ECRAkWcNiEgq1OznmaOlFcPm5FCe1FSj7z6BfshoW3E8i+3UfTROGAO/
Pz9e6Msf1kZEds5xrGGw9eYHabCP+tHbp5E4S5ZmSbN2PbLK52DpAuUFhv2F0K7vbj9XwKMA8WPl
W8ROwvMl7/wqLB3nXlLcs8Ml6sMu3C+X3fiKzGD/re0ubJrslUfGvtgdZHuPwcamqxKVmqb0NYLT
a2vSg7dv8ZMvUwBjXW4K4vMgp5H62ILJBOb+QcIuYMGHln/gVPBS9WlnnQ+4G5X4K7ffx6VNIpMw
jfS+Q2B5vmz7zp1InUdZn7uZFh5EJkOMGpj+MOdgBLrIdncIQi0xskC2zD1Xm4IJ4NK5lqch+hmq
dvY/G8ie6u4fj481ctfH4jHgFh4+l6viBR2hI5sa/ye4IMtsT+gDW/QJb86qjV++P21RQsSUyzF3
RZkil3GghpOZs/JD84mhBdbSDabGI8eF01JEnEOhWksepd7qWM1HkXPcchVyx7yosT7begl9hs9V
nsUEdklnUu8IH5QGgnmfjA6D/q1OlGUoQTXL/NaziQYJkjSQ7vAQOz+jnhIkaSt8Zabgy4q24D6m
F9U4BkMUxG83Oxp6bqn57HCKg3rtyCTDK2tl/Dgf+Thyg2ajOk6klLFvPOX7VUxevp8mPWfzVwAL
qHHh/XatfRe5Mlut8dvL8IX7yMjf8QDwft110CAezfr6gW7XpuypQNOvyHwuDhDHAfdoO60t4Jlo
Yt5vuh4GmDCZN3iY/V3XiMpWdYkZIMqrbe1VUwuV7/RmHnCtCYTE7VfkBxY+RFiA3d/3O3V+7Svq
BZxnZJeQhGncKns2nZZX6PeSHeFoq+tA18JJV1khio4c+2isfSUTzP8jPjgM8Z3cKqFjXQPuPBkt
4oZgiotQLiW3/dUw5Z9kRIrl53jilQ1SAoclNOvcETIfyTXtCuagix51NWkBIDljlatCgoHMofaS
p1Ag2tZBeeqPkz9C4GPXlTwkVaOrFseXUvdrX3Kczy5+fVUHISl5NbcOgH6YAZMOnHdW1Cy5xg1A
XRq1wSzCeCfTx3dbhepj1xpIwF0mFXopVSVm9aHkXusrQrJEd+Mx0jKnv9iM3YGmmEXO9Z3l94aH
pmzzAmD8X2poo3IeTSXNHj0Cmd/DQLuQ7d6cxFzsTBpXo1SA3MhQa3bsFnKgqG17ZPBe3k72Xviw
yDva9dslq9kXE8W3LK91eSZtEgyOwg8unsUKkB/Kz57p8i3iHhufKMKHALHJ/Q6EeSt/9zpl1+7p
1B6rxA+imCJPb67rDOQ+vU4vWsI4z9tav/CXkyEnJNFRUHMxx5gqpEn4cWSFMzbq37XQ5Yooo8lB
3g3TmKtaqDo3Em3tx1wQhzXYV+xq334xlh9CwX5Bx13yvgklz0nmO55E19gYT9bfj9nxNt/ap7RH
HXAU4LO5H94/glVc0Kc4XZl1i1GEKcFhtCHX+F3QulzuyKv+6Y+OgHMgsT0kkbAgSXOf6NcnWgnB
wUJb+KlozTNHuzPtkktoLfYkUh9T679n8EgsvRm81f+z1f+EpsNQBUeP8UlrjW63LoXEA89lNRmn
+0OmndXPo7OTAOudfbSsscw+2nIvy+k5n6vhL5x4x9heaTTlsluYq8i9BbYKT3FdQhirFdpHSCsV
Jg6J01MMwc7AV0tkL0zpKz4rtJ8KAklPPrWPkwNS3p1VLmjwWwv6BNB6UvI9EW3QDQoDWVqfFG93
D52mecs/KawglTguwq2MGbl8VE/tE3H+k+YBjP7c3MDblATZG0gOmQT3kmUbDGe5tQp8PWHvRPoK
cqTQvEY6CNPMB8Ct0fAgNcMocNKcxNTspUk+urZR5mhDb3Fvp4zPGuo9poUyg/K04RcEe7D0GSjt
BjL5g330ePcsbNd3vGdzPGaCy0kh1RYcxx6uRt7Q7Cw1vXN8ESh5Np9XuafLPksPqcNOg23IIPpY
gjypzr3EypY8uAH4oZtX30+a0uroK90i2Z2FkXIUIzqCftoszZiSksVNJGcMRpOnrmqK7P+06hcd
UG190UVOer7wz7B0BXRkKik2Jd/0NObX7669R1N53I0SJ9QYjkYPlt9ibZ07mbru/mpCel4yrnHD
/exw7WVJ9c5WQ8OTPgbsC6FiQKUYApz9Jt4pnqG6fM4mKEq3DO3ONQL2RhzBrDa3KZOA9BusbX07
dAqSu2Uz9XT/jKTQoeZmDsJyZkBAFWBc7BjCwM74Xq9vctxoURWVlMiIt8XOEyJh7mXLF3Ttz4f2
G+cl8D7wWn/tIy4guOe6amHM84nT/aRR9UIDk1S2ooxKR/McpAHnGti13pjw8CRvpNzRkeEHJL6K
V5w5GLBgfqwDOe0STi3P0rtiAjqNFhiBekNSC+g1Vx5VA9LSVMJDX3paPltH6r+ondCvP953gfvZ
6A/ufAusjGHbuJm8ghkHwnNQPMsUy0NTT8UTB1LMD2kuoiAkRX7ij2HuOdFdFAD45yK4mGeqEZC0
fIICTKyc9+WWzFDs0Bf1hGEC0cAQeUXzlBlKkX9XlQzBI6tdN/cwLmBRW4GmXCTyFjhEvDBOmwmj
YtO5UQwHxRFtrCrRPr4DYf8gW0F7ZL23hD2L25oTqsyFnCRbWNvEgCpfQg0RfDY94e3M0wUYYxvE
+5oMG8uIkAqZNpumkimGmTWKL1ftod/iA8KARJ+FQnVHPeHdavzKHWbD/St9soHtDGzQhTUFJo6i
dbpdvvxKZu2UoWOM5EYck7p8xY+kefcRXf/pBTaZ+hApLiA0kQDmf7dACm2l9vavkFmYuX3YeQS8
GkFgnMMzwxKYog5Di/pIbUFT4728nFfMfZkFYjO2sOt7vo2UCG/qxu1EYz6dGrIayBDrZUcGx0So
rVae7sUnYwwujWwlBd4mtz4TksB94As8xz9YTrW/7gdTiXnz6H0wHHzFIPxMUGxJrSvr0owDGmiz
970Pwsg/GXFDdqYYoh1QQ5fppAUS3nrZlEGy3hk45Qj33Y3aLFZaUve12NRZceHGH8InZxkdz9om
9xoeooSRJ+NtIURVft/9YWsXpABjUTcieDTSLXzP60C8riYhAfnhBI84c3LsXQSFgLMX1lCm30Md
p5rmalHUsxBX/2G2j2e/B7ZkTbK0dquD20f9ObFEnaqsWddElp3VTgO2pLaUeOP0rqm2G7nrpY2j
9JosJYuUbtp5AXgmHmA7uRSAulNCnDmA1jVZJoM5n7CDjI6E3EEbFJGupNv0vkjQ/zh37wvd6ezf
hjmMVRUsA3cQqZLAjC22r59OmnNXS6D11h/Lt+gt1+cITk4DZISehB+C6dfmD4QSUsm8Acf34OU4
9VNtcDHICgfvhgNr4LpzpALMITDV33WvrIWtC4vDIHtI5eotNdnOUI3ppCFA7EOtXnDQC/4ebSuC
k2NPjO3W7HoLupMDsaPhYbp4Bz4NK8NjgNZecn25pCIN7RKTwVCo6o0latTKA24qGqdAok15hH6o
V9bnlSseGj+Rp/wVD/AzljY07pnm83cScCnBWjWmHYMOYfMa+AzSJkJZnbVV67NuQGl8/VIeczdK
99Emq4i1hQNPExmmpIkyZ3gjSfT9GMkXZ9xtPDIcStemip8nH0mWL6+i40QIvkdcEL3ATVy6ti/F
UFii4VNEIyrlpGZok3f4FJONRbGGSPhLdm3hpNLt4keWu1R5bnmpnumoL5EmhYl/TTE6wzvkHIjk
eahKLNOC7UFPs6zPIa90WuVCgMK3TXXFX1j7MONse7jIkH5gKuZcrYpY5CfFz2qfPP14rm5Q90rp
VzVlv5aTe8fDHWhH4s6/eFed/wum5WS2TDhp7b0aGSOYuVMt1wqwB5rfkgAjx3dhdLrawhJ2l/Jb
C6Rl7dJb+8i0lyyzS2pbELGXLnfNzfVvoDSmXU1XlSEcAu/GcG6v4pvNz18JKH5V0SeDjXH1lY97
kAw/gU7IpLfDyI+4VJUfpyoEEx+ggDRwB2W2iHXX+wjBEP2wJrGyim6IJ1nZORMFbgO2IozWPkyt
FCz+C4jqjVlWaXJR9QaNgm9PEC1oGNms/P8fJ6YXuCRqnFKf8rAem/ae6fq166lzx4AC2BQiAWIy
e1rmPud/hMOdcZ2xcG49F+kGy2nVBhCs7KHyWEN8bB2alizFdR0d2KeBJvtI2sN4x5bOTfsQwVIS
2itidlwyfJqW7gb24qaaH4VCUUzaLb07en4sGaLoP/oDk05ktIGpfry5PvDSHnDpyvBYXpk80YgK
7W5LK/aphvWAeJTKbkp9Zo0AS32pwzAtD1PGi8TH3gad4BpW/xb3Zid7xuWLskDsCzoJfL6mBH8U
+l8Ut5Iyilv5FY1sc9rRzFZVSslLijCif0VMv0+zeu1S3Is+rRhTrd/0hLcGnQVcEWQYVTxtSuHb
gs8kLvZDdvrhbCcN817TQFGXhlfmLNdtXKMDhyRMQw5l06w870RG9y4qctopVmY+kpT0XbKyZcgi
09vVpWNlg5p648jMAsbnEf8dtPyFTNnnhVm8buJAjLhhdghmneJ31fLcipNhwDBSqolWdsSQUTK2
+Mm85ZAJQenr8mEJiWxhweyc8xik6BvVVW75n0sphJzDuXbHd2FZNYX/UjO+mXGcehCzeS3JEg8+
3clUM+eKsDsRncYuyib08pnibD7/RWa3Fu1Ji3spxL+k5sdfcSaMQX7zUkZRgDoGUKV3hU+/aHCY
Q0f5EmWhUXss2s6aLaA+WMPY0iF6LAsPpqKOcDSGItolnVqIo9RiR8Thgw7fjl4ieJ1hqiULL40Q
WUqSU7xppTSmuJQ2zd5r+aRNyojtfKI6ZlRGYJKENgt/WjA8ONVe5zi+d7Tx9k/Me59OxTmHSIyU
A4/VqbSyML34EXIZqzwoqcDD/WthXg2nIn0LrU7NVYMQsaTngtyzclPRXAHlUmzrvK/hNLOZAtxf
79Y5J7HV0LKv6T+tIfM2F29eY/hVQYyJ1Mu2JiXTcvr+1DvE3sdYYUvWnu5bmIbUh45zMqArtDrp
iCDrwvtaAQoAuk7Mh9qUGbOwnzWparcnjp0AE0Jfdu0WRZIOiFGfBNSffkD5wYMQgHvo/H+lwbF9
TFAKketXo3cUKpbE2z+sABY+3JyEL19uFB8iPEp5HP3g9k2hlrEEzZb2pr3qjBxpTc0wS2RPubdf
ZPwcilTfMB4nG5dQdLGraRWHIaWSvBLylxonjKiAxpA8vB1QtT2sOR4kCEIsZJtFvSEmaZdi6AHe
UiHZykSeD1TXDQBHI3pLJsTRVfV4gLOMpWhMjHh7u3hXN4ti8njID5l+kLcjpVT0f4qWxlIDFTea
TUC80jlSbty7reiTdqSKilGteBdl5YQeoVi3mlWsD8SR/hJ7mj7BCZ4/4slBuvxdChQAmFDsdwdI
g1+DWvTy+4b1dmasxqDP8eLpv5M8QoFyhZpNYy+1U0yC6ZGI/5ZpCdY+ZqctKRnj0PmQGz7lnBCq
K4wXd1OfkyTfgeIP0qbnlMomLl9I185AAF44sHWXoQHDY4TrlhoibKkMoMpovgaAQQKdr3l6ez3W
TVB/vKEmb7CQQyiAx2cW99XTuWzsDU/4V89D2Y2nKeNP68e8lRsN1u6BYLvRM46sgJ5s70p6DQp3
CDcsUs1lJxTGZe88eUf1yDxHBrraFJQudngPQ+93tyO34+0HsUqjpeeLaNh2evfld3l/EWPz61nA
RAScHkZ/O1t1UQz21vQAHAlNiX7syqG88owImfYS4jGQBw7Hr0d73Mh1UMCES2GjEoxlhNxUB9er
fNRBuUZhwuMKT24aJqov3H6bOGxcp2yaAul6gxRa00ieI2FjAxy6L0dXakBb0eL2tsMggF1r7G6f
SQFIrnC7tS0zaM0lOG1WdotJ29nFaawy5NjB6ZIPBqmykavlfuMb8rD14cWoTQW0nZ0GZC4wR/wW
BrplU16bMNPhJfitWafz7bCln8YiLfv4i44T9JMZpEt67Kims5KcDLT2nz3hlJ15i+nfOu3im6tD
nD/jmt9ghTorW8HGaor4EluoCiBVXLTfyassIa2dchqE90kdypLJFcJz3NJcxXMv29SYBQNI+EFh
E8pCrbgmxzCAH7qlzQxD0XrT5x95TABnPiKYd5R9z0pSaHLHbB4Zck9U9yDxMIVlrhFVlY4q4+rg
5OZ2iDJ8BHQlxThJy5oF2yU+EH7GCKP1Ab3FoaEa/B2vVMN3ZPnjWUH7Ew8KodqvP+ykrbUcsbXN
yUanNhBj3FqgAMIQRHSSUiO6aPLyRKHxXkJX6xHdok2DIE5F5Q6It2kCSRZs9L9e0r/Jw3/l3jOG
L1Y8eO2bbUCwuY/YHrQw5IO8vi4GRwL4DRT0y79SfeqfjJk7nI11fLyoXU5yis9donfgW0PxHWtd
UTjh4xvaikE1HCoSWfPOJMIWTapqBcdb5aModHJ9cS986OSWKnHJ3vN/ukvbsIE6WQzmHhN4bwpj
dUh4rkPMjRhk+a/T0DlhdR51g6MbGXaVCzBCttcww5nw9qsGEzvrIGLV/hvdaVfO4T06xJ4xQiFU
yjhHup6OgC17yhytZpUFGkFMNHQ4qMd1d+eyY0HN7rG7LvRDdiF8LnsSz9C8FOB2BN4AFxKR0JV7
HMOGtuOLG23kTR8B/b7Rosd+VWX7XlMgfPO4YiWUp7uNIiYD2bJQWcDfjzAm/6Ezt4xHuxOGB1uC
YyCOc2ezHIqT8FP0tw/Waw2hyXFwD67mtVQMIH5+zLm9eVlel4tyBczRflclz2HYFtl1zj1LDOZn
XNueWrhKnZCqi5Jy2C7nEvyg9YWD5vypbef68zEMF6OPxadzZDISRcUwozcpgDNjeqqPcXiLVZQy
Gquf5y7aEuu3zWRRHG8z9zvML4H2dHYC+jw68C6v4PwadsK+idBUdtir5DKqAi72XLugi6xqxm8S
LOI0KPDiZCttH1OoChTHxckakjYgvP1tdseBs7L3zMGnjULh7RflO9k9qdPHvKLkHWfKkR9pMbBr
R/vStUKAw+rNr6KTcpajUxq9Zy1HGSBESEBRXDwFC3UQLk1/mRDT/TmGq21uSQ18dBMSgl9l7LFF
dhVO7clY1WUKkirCmZoFKlCV2GvTdsQgQ43lY7DrtsfQW7eQpu5SXCzZnlV+O9iDMTqAtuS8h4RA
REB5aUKqh7xrzT8oOZXoajLLncU6nXk+8FT0IVdKXFZ99K4E3ZRG/LUH487dXDf7SJTUbMd/FJ44
pxTOfC2vazhCcYrBWHceNAftaThpu9AdM+w4az7gN6cdn1V8S76zQ8zIBfWDGCrgq9j2IZ17fyqW
uJPx2EN0PVyvh5c0yHpoNtPXp16cYCdTFaWo7AgA/PNSlXETVscfoxpAAYHBkJ/31HmhCzNgIIJ5
GhUomTU8fj4HAPTQnkogAgMy260D51MRGrDW4T6sbIKyFs65golNVLc3/L13M9a/rJH4PBcUE3kp
fhuP3BBW17LrVJeA6C3A34f1MEgvHJvOqMijMuzBNCZWbJBCzgh1HorB5V4vU6HhosaOHv0ZWf8w
abXUxa6cSrLSstjjXdVoLv+NAmCKGun4iHE4gLo1rPW2IQ1sQgNx2Zcxm8ULmbOijoPEzPknpAMI
q0aZAfuLRGw+UkAuShgHOZTWi5CV3SEserqE+1Cby+LNksrTxitLKwGW8HRqx8TcqDjTffkNGWtS
xYfnIdvFYqed+6iPllG21YZR89QLzHT5PPcaxSmJjJic2kVQJuk85tihHngGI/knUq8d2hZQWddz
gg1Do5wapp2wwoTW2Da/BCm20pDbbozEqQs1nZjCdS7e9L07BEWxWXFIe0r89JpnlGQxQwMoymeN
75hp3svMy0iXrZVy0nAKLk2nlX8e0Urtv8BpWZY5W363xaDLT4rHJJ/Wxv+SzwQBaiEkahBws1Lo
Gx7ii7/mdzZd12Jr5TFfUXoIsu67EJmHKp4vFE2PV2gkjIL7vQBK1kRAC5QJ9V+C9r1AabCB1mvI
9T6I1pkpXuDfUYmkzLMpH3IP6tniQBEVWAvHNQKTuczX4kpqk1XIUYVAe7FNSIMGtN/BRkGSsfQ1
5I2oBS6BCPtOT74BeTAGAT2IlsIMwe7PI4T3PFJ2pR2V//5+gplrV0SmSEv7YRCQ68mu3guGCZgO
M2W8HBI3g7wHORDQCX1SlyGK8wEd/712ZfBcX1Hy/pgwOAsNLePWoeq4RvL0llyD2FFq2C1V6toN
wQDLlcTCcULdO3hQmgpN5Dd+Q7JoF5or2iPsSPl/EQM0WqnDHhFitPZ8IZ9G3ZpJ8/wWDKhIWuWH
GH7nQT5vRlFINn3rtDjkhJmQLPl5Zv1s3jT3UMd+sd2cpTtopqevGrbDN5ZCKlxNhKXPtD6wr+Lr
22gGe6T0bO8dSHGLyv+4CfAakDXRaThP2HaHIAD7ZklPZJXPNdkcTIHe6q16RO03TH6HO/J8767J
J1aqBMRqM4AbNhR3NFzsOZyP6QpyxRLcG3PoCAhK0w2iC3Agiyfben8+47RmvecgAT9dGyN78rQ/
EoGLHd0lFhTr9xbsYRVotySkSc9/2usaD5gxRJBS0jEeg9ObS/HFvMGB0oJklqAcL7DUwv8VOHYj
B3hnur0VK2xEbklQNrlzfXZDu40cfSkXwD/yi5VfldhklkJH1xXl5/7V8QGJhjWcV9EnYN1SzHwx
Qykc0df/av03WsUTRSEf3k3Vn9nhOa3UnRAlabjQiPJvUskY+RFPeuEOXe5WCmEfGShznrZKO200
Oxvd2r/UbCymkKv0M9woivVHMo1+/8POwR8tOXRVzxKQllig9lUnbJPitybgSTOmfypogJ5lUw1L
v/8DrhDhXaCUoeVwVU++8ZV2PHpzgdb9uDe5u3DiKzFsNzh6mqsMI8KuI8uHnTlAU+Xq4yZfnu8i
l+3oc0mh2nR8+wUSsRL9XMyMZiwLuvJb29KTZRbnP7ekUdk08KA3Bpw3dMflLY1apr4vRpGzx6vy
J2oIo8mRBVv4gB9jI9sqtYcgaRFvTV6TZSLM4UIdDlyeOyU9Se9oOaT1bKZxP/epIhr+y/uQcq/K
jWr9JmNdadxEQEYZtGlRSYTVSbJybTp0cX6BtLv3W524Pd4lukl3Jo0KTP7hGnP6BgK5a8JJlscT
v9uQvEAqdSBKtgqhuSYI61ZD2kajU9SlZG0cDQ9jzYBPxDt5r4gIPlwRcElMd7S7oOnP2DaGVYzA
TAX5yOpJBV5yJvH/EoEboKZ4+Rve8/nyszwlEEDAyDcgqnnmW+If4K8SkDJ2mOOheMSdIHTgxqBh
On2rBfrvZVOyiqj072ihdvxkdv8k9dA1YDiROhgYOTlgdbjZ/gk732fCd5XrZtStZN24/aKZtOri
LiVco8gb+M0TiCNS8MWYH7j8h5zl8NlUAEUjfhsWdjLywiA2KaPG+LMdf5sjOBuk4jx/1GOOQRFo
RkCtpJfvtoxsFg/YNA8R1JrcbbvES+ksv6o18Y414pouT+pa2p5W9vKyBkdYsUAN2Y4WXX97PkHO
/qNqiIx38qv6G3XpS+6zG5Rjl8kK0bv2tPRbu6ljqQGd8BaRukak60CvRyK5DU3b7i0APYH+Mni3
ZPuxStgybOWKA5gVTqmZYy5Pi+eN8xPhfDqt/vr6wofZONanDPTeg+z3R/XXafQE7RmuYe87k8GC
w+r4I11d8X6us0QRaG9UIMaWPle0D0q8GZZMyDZrUSO0YA6iiGokmZciikzKHdyH9X5ub7YpXQqY
+ikzijOozqn/Z9l4C8QnKIt2jbzv9ByiikgZ0m727ItNTBcSwJdU6yafk5um/RJrieV/QCuu1mDt
uq4/KWCF27em3ZwfuKoMMI4XlR0eNuIrJ/wDZrNTH7LwpTg1Kcq3i7FieoCCX2OQmMPSYs5Kjicq
OrbmUHuwor3XuKfcbU90IFP5yz+nXbm2/mMLWlqDCus/UWsU+WXPtBbYf0JhkDjrj60Me+q8KPLu
NJzzRTj/36upZYjHa4M+k9L6dF92MxktqIGdGaSZRUSw8xFqNqC0H6TiIyGz0QHSdPYKGVcn3dVI
eyV/PlfbhLBAAIKZby7t+LioE/kYQli/mpmq1o8ffscIOufwLLjfBFWs0SNKsXEgwjaohM7Yx5Xo
/yyE3Xy+iLFzKvrS9ERkm6uBWOzdx5ek7FOZpkThQFtK975SNenqjNUI3r+1ITHvyMdg2mTYMmV0
81vH6xxSPgQnVitlMrIJ7/cnQERn8rgJXMgkpvxb5zEqcdRJV2jv1pEjd6bE2S78ASqoznkc2kE7
dSukDlUJQQ3eUEQxbSOvcqN7x8PAoCm6ZHKjpsLrJVpe9qMpZujSSkRRvS58PBhSzG4O18FAPyHm
u+puAk+l8XYewvzuSVZJR3Pt0aTk6UqxuaLntToC7uLZup9HNrfBz/ZGjVoJZVAZbKXhfd6Xzgjr
dZgx6tQl5f6kXI/Tpg0PvEKa4GUYNFkGW2gNDAjjwZfcRdJINzzYJiec4pnN2Xf5jVDCUKEMLBwm
HHPFcIQa++TL7dAQY9pkedoCDevghfgr4i6Q/t7MDcbUDlVBSY2UW+CTKXv5LxRxB2I3H9YV3h5p
bejhbBAfNhsWZbwhzDdvnWb5y1YjdkVqLXfuovysm7lZz0B9FaXBVedcI7qvhUoLwkukCWIMS/3M
x1RWXfo5MaW2fY2KIVzGpEgWtFNiQHyTbjb3EtlfscVvdyfYKOjCdQ+9R6oFXVAGADKFDR/8fZvC
BdUjwOb2WehzuNpBwWTIIeyyO5LReu04lnzxe6Cr0gdqzKqk3gsdqvcGvn+Gxfgt0q1ztiGZQVc+
XA2iOFSopeDoZrlZkhXJDJO070VExntHDWilIZwNZFuAoUQMxYCBSqRkSaG+AdZVsFXn2IbZiWkL
m++Pn1wvb84bBykxU7y6khLTpjJu4WE1Bc7H3KAim5VQu3YoU4vxXr6ZdOEOlkNwZpZqIClLfxQo
OEQVjVxJ7HO/nuYWZi2JSLemdVrD3lh/r/jaKkhswPDO3onOKBPibncUuFBXR+pK1a0AqTdu+d6r
BN5mybQrGu4fc3DOBcLnOZZ0x+m/ro65xdZsRWd86q21hivDdghq7dkWNUCR8bHCNxlPevxi65CX
QgWho3R3FevQDvRySRejw5zQhpdDeyd/ZFnX9kbKO76m847spVlifCKQ4kEAZckyFvsFXslJ1Zvc
T/Pg2JbILPp8xsJno99jH5ZCfjGpelUuDCY/KEnLbY93EFuRpHPY655loa54ol/sE9bDhNJpHWJq
2/AImHsh5VT3HKopMN47DoaNy4OvQMYipUCYiRuk8i/g8WHyIlRlFx0yAEQKpX9hb0m10Sno1513
Y4JdZbdQXJ3AM9h9WMApDLOcFplpP66clGzm4zJdy1i1I9drmpC/OUwygOTrK4RV707q4QOSNzZy
so6YClEqcVpRp/5M+3ocAgRo3+W4yck/1m/lxa+wCan6iGGqTPm+3dfzjW/QFFiFE6gzCV/X833P
LpM1siRu4Ip0W5rVOnS8hC+EfICCF7r9OrxBjKJTwO3VRB/AXpSfrXmMOCgfMUnylBVeJvZM5AAF
32WinjmwBXkZbaJ9yqekHstltjvga0nBzqPOzNBES/blr2n76z4gXqnUTX9i+1AruI76Pne91tsl
IdNpcMdgytE9EY9svAm+VfFY463JlHVJq+RBS/k+XFsiYB0R3qOCX6jU0oO+SWgHfVgITbMfYuY5
Hj30sx070R0PMEQxjo3g790SX+cTa+m7+mQESHH1mlKKnN9dgd45THwqxk/6XNaebqi4Tcj0hdiQ
7cj06Un+2kopZoI9606AN+cHhsD3EZcZBgMDiuTe5NdCiyeXhEi+2yaot2+i9+IMJUY+uZKKAVdj
NTc7Qv8VsGzRK+uAjKPMfI2hx2nZHtJEogw8iRjwaLYB8o+Om92fmLqLo96jELdYievTQgAXCoj3
CdIjBxSjCNnVNtW+8leBywsmLyId0EYi/FIQfsrtJ14brQkfllLInn4XzIDpWhSjtWJn/acC84Bu
8L+Aqe563CapFzeeAYQeHOAfYEABHNvwRpVsiP0HSgfcVogTTBdJNI1uvyej53kQSEiNOEprwWIs
pFtK1W/Y37nMT7dZQbYqzNBITTPtdZbj4PYC+wCZ0/k6Etu1GMeZIZxetDlLZzTczokLwXSggpkE
EfJBRXCuivyISWacaANNP0jSYX6fIsSrF1yfLzElXXZlFNNmQwEmFHI9HvtQ1LyiytS4NETgZChh
eyXk7GrHvE55uBFcueQ+AtovR95uGGJTRRUHo5RYQMbj7s/Rxo3ldSN1u+SDRdm/M2XjS8cmHa/r
iUHTClb1dVM4+S/ndwI8RKw52wQu3fztyU4PrZ//FbE6ZLZWA1SDITfY7bH1SIYIw2IGeX/Pj4B1
DpPQmRZCCs0hyhPy1BTkLvprCt3Qf1SMOn2QgBdUx9AAUZFqXQwvyv97DkXH2QC2TpJy6B+qCbG4
AHyDGnLwpeP1D42p3lQGN/X+Pa3IikudGE8ddpqEomJolJlL3nyOb8UWeXY1MBhp6jkDyBIFSY+d
YwWQsxuee3UWOm7vHb3RAoO9PxIYhAJOIbC/aRR1xNAIyrHmjTBI9gl3kZnhEj40jlhgEHMVdcgz
k4iaDPWVa8C9u8qeWyUxuV3gTnOdM1TSPp/RiT80Q2m5l75KzgM3gv0ePAyUhn4nqDJ8hftKUEKk
qkgt4Y8Gp11nHwiO0Sew4GRWsEvNR/o9pRFCN6pcytp4XCox+M719rSsnnIYUkwpu1gGRq+3Mm5a
7wXaNrNcqruNQwR4Ny6mVTd1v4fJhHvsNSHTVW/ldtoJ2/CshrZwxewAueoLA6so8AGRMHaneBZG
KxO77icX6H2z2LeX43EMtvXqegos0VRCWlTWjmyZ7oDO13fNwyYChesdhM0y98B+dvKoy6KDO4Vw
O4lfZ3iiV6mBMIToYS+saHC2LxSbV2V43s5NKPqbH0/luV7/eqMpSQgbjTuuiLt9fCWXZEjmGJnI
Ttj8zAbwL4WYDK7NwE1ngP6wqHWuQOl0BsyCzBP1aUrvyA55S+gwr0RGDV1P0IIPnVFEHZ+EFyK5
dOVKL3WdS6YhYKFHBX2TJ7HONtfpQlM2KvGRZkYTAyt79R7R506tagAn/1D4gGIXy7OvShFM0gF3
N2Cmz2dRDb9ptWveoWCpNTGqjq3yWR3vlHR3eD731a5qNDKQvrQNqH4yjwmLOM8a29brSLLUOCa0
4+9oHj15QwUBwvj2eUbplbSyNnCIARPDdn274ZgPvu/RtTylzY8UHLt42hOr7x48rjcnza9QvNbU
opihmvf+HdSWm5KwL9DYxK8LXdv4+p/lmOyqd4yQP98xrquJVMOPmWL/wA6ZzyzZIESCIBEgh2t5
VeDstNUuOd63A0k0WR1r6Inwn6YraGRTR9SDf26LyKOu8TmPKYYDWCt8g1Kozamlg5yL6DR2Kt9X
nrrn9xXJazdRdq4fyV+vZFpsqaFoQ5oKSkw9IHSr8D+VTGsSb55zbZ4gkcWPoxqxucNI0gqo5BMc
EFscDclQ/zSC2Wh5mjIdSRkhJXSnv+v/0ZRdI+zNtuFojWCHXiiNZUtw+S7rms7GMiokDD0YvZqE
o1u7BqMAbjmr/N7xvFrJhgiCojSFBOslGrPqiE+h7Zx3eNncC6zcaqgpXHrYcuS7GyRa3mhwdxaS
ukTDJWNL4HmCKas3arsXgR/nm9GAIkct2OuND/rcrO/eqCN8PniOv89Gc5rWZggQN48OYWNznb3M
aZV3awAYgp2YZnCX9DVMIOzn5+M6XOHiGupsQD4U6jcpwGiAuhP2JP4EtsoeBLk1dU0sPya3kBRu
3RH2h/852m9m+rDcvE1a4SWzoh/A3rTu4bMRDAabL02ZribEOpkoHs2FpgTL3AWIkbrbHb2hD/AW
6t7IBh0iOcZCF6GY5axtAzNXyc70vCRN4HnO/H09VMVein87dTP17puARSSVCHetNzwEYrrvxU/e
IyMJVcMMnqt2EIwMNSMQl2yRh5P2n+F5eKD005PmfiNVutuQBMhbZnR8hBNw8sTImIyh7kEO/8bj
cH77A/wHpbPhMbK+LNk34ZkztoEMN2r8z+tL5YKmKo+Bd3EEGf43f+G/pCHqR0OzsDlPvXoiBivD
WRmOs+Ln5J8Go5/jE3tLImifwWzRb1lxE8WtkubE56LuCJesCyi6EZcEsJbmVtuUnxLCnxD77guO
nKK5L/YTu5bMhKAtLS+JLa6z2KLjjZf+3rcDEAEtgk8LCkCCT8K/KY/EJBGKyLa7dzeq022XeKZ1
ITPf0imu77kNdER+lAoyMcYA0OYtyHNgw4zPqCruMfKJIBnUC9AC83mIjYvcRzs0O7qbqevPguKd
Ym1lKL+bHDZhrgyA5Sj8y2Dd5GUK3aPA7DMDyuXS0kl232c8523eDr/HmfVLaPsd1JNoe/eglUCx
9NfOVEMmX8JG8o8PLGcTG9cPvuVZttb2US7cZecaLW1Kq/ld2UlhPOwV9+RcrtFJqKkYP0x+NNiW
X5DVoZeTk9OhSLWbvj/IXJ3VC+O3TZ18GbDls6Tr7bJ+YguM+cs1dJK7aswQYcBrpn69sqoqX3rJ
LngquyMDiTV6qswaK+w9aqGrBTHpZMiSIx0Ou6UW/4+oSlzmPfA1BtVIENPXi4ElU//QPBQjkB2F
Q2C6iA99MXlVhyTovW2HCsSC9vIXw2zgBXrpGwGhlayfiStl0v67DKEggkbCrNlIfht+VEoJMYw7
kDFunDPIRMkeuNannnuc/folkrkn6gOaE/jlYU08YRGHHEF9B1uPDRHswZCEpN8YgT89d7TcQy8d
RWLoRLQ7Ey1qTyL3/+jL0zAGR6KutmVmlLfCm+WZmE0J+Tz9PmgXSPkGHgm2czvut34/9eAoQx07
peuwkt0BulnaCEictLwYzVlisPVcUdPo1UDqCIV5RsjNFiLkCa/InTYguli+SHdlmC/nBDb8FX0F
u1h6dJy//6cO5SAjVHydbHLQl3o53hYcVi2b0KNIS9gGjjdUie6+Cs26kOYp6GhSd0633CAf7RGS
lHoViMiSgXt32fEfMNU60PC+7I4NGz4xEWHQ39x+sDlGFQmZZcviQB4K9OiwZMMIsTiD4qV/zDL1
Xj/1lrzYl40XxtjOhn11/tUabmbPIKKKgw90W78C1hWCVoOEV3rL8eHsb+Z45v/D7snahZPjZlx8
sccyIaqUfsaXorVLkvl4DdOAwta4MV5ITJgHg15/i1cf2kss7tJgrFzAJ544MEjj4E6WYNAerc8T
qLPqz7wat+E8tXhv6DE9X+gKZxmaghRh9YLiqMTHV1eEsAHdtJ9jtFRYSNELZg7W9yBmPZCxZmPn
XdIBaFn+YOXRBVUWc3RsNdBZHjL+1XnJChGcgN+N9221mah3PY1pW3cFCZTWGkV6lFqHKw7PyIfF
Aa63D1As5WchnBL9DN9s1UGQd5n9vKKNgOAAZMCcK3bk+7o9UAMJ3IOsI6/crlGUaojR8SkN3Dco
zOKhDPRCo+Lb/xKI9CIh9lZt20VanERaU1tvp8Z6se30I6+2zPf8ml6u19FxlcUmfRgT04WlaVS0
EPQi/iTUkO4Nn9nz/lCNXbTIOx1SzfqLbWyknMtFT/+e7L6FbGTJo62CIcANURNO1bpGWoWXjuj9
hdnsWxdNp5c7sVgNcKHR+KMsDJ3fk/s/xtcwzymbVaAP/X/7K4e7uVVRKaPN+U9bsYywefU8bIJJ
FQJ0PZnAnROD7rImiN9R/k0Nh9ZAJxNfD3fHMKeegxgM1KxRwwoIGkF5ciLIswr/DuOOeayF5QkR
fZ2kE3mKuB8VzPhTrJVAIsUWLWOyStb/iFdnWHO0FFfE3eR0TQZ+PFNAhgQYwFB1azzUbFPntGIH
xfEQfmuXRPxS0mlK19W6ZKdRzTcaBOSzqnghm8HQ18lRRLiHhsiKXaVayjSmbsYPFGebxKUA+N0S
GKEIt3KhP6vipqZvJuLdWBZYNBL7tRus2a1aNjD17DHU+5w/TI5N6g1dtS28s/JqTX9SIp8k9twX
GHZVibe92kGgQki2CoywW7usCu4a5ezujM2QpjB34FHH1NB3uj0KW1cFq3Drc3W75jfEj5JDPiXA
p+l2AmIlhwPqk5bYx7jnwxbAxXOlS2U2SIXrxJjPLBNw5d7hyoU4Btj7SQlZRXVb4buR0CdSGVxd
IvOryrbFlOd1ZJInf0TTOtfZ1gMV5+cuvKZAISNlVdORkmuN0QJyYxBpgE0VwWHG2oAGdDAcgn5u
lJ5EiOqlTR/IR1w6NrS6D+2hycvYmIIMpyXtWvN+wAdfR5kl+JEckBdOiizhDnZhzIX78zl21lsw
023rNorK7NzySqFSZ82Q9sriGlBh67HqTWPZaFlPf5mG/0mJL9zni13x048s8zcaX+u/J6GZDTJk
5Rr5j1c+QWYf1pkU2Uj9cYOZaxFzDcXcfmZ0S4bx/+Jda7uYpEEErIb28Yy3HHiwzcCURfO96gzm
VvtQKYP0wh9mWfRxhyOjNbuxDywB067/7IoiEQGo0KigQf8m/houMRL6bpr5gfUZnrC7BZoADH86
lHi5vzM5tDpR5cR6iCojJ8aewjxCti240uyItLNQQ3qbhrVq2eXusNf9nmg47ugbDdHHQFTuZCpO
dIgNY9bF2BOzvgPxXyaokKBOY8Szyr/34FuJt087AwAGT0ajw/9za52l3kYWUu3uZHQT59z8Mf5n
WUCIDXCb3dPUOKUU5nTAkp9plpdJDMgY7ln8HhBl2v+wxgHrEFZNMdeUECskSndgdlRpNTRmcJ/1
rRG96BAJLF3gO41nLsOZn1ByV2IQrfLKXgbERI1DHoHMzEtJnFHnHTKNjkaCPtb37qJnOusHxe4W
D5tWPqnsLQveGZyCi03Te7Abvtcvy5dJOjgwb3VzfOvbTKkcgcurb3lztFoLjefdy/ZQsyEHEJMG
4ZqBGNhILbTCg3g0v+bADYZFf7U/qE4hDi+KWxXVdgsQuOdqZWThDgwiU3XRu3jYO2RRcoAxNpyC
EX/SYPnvFCZg3k+M7L1vXO8/ty5TO2nwyCujAdEECP7nrltVXjuyBJBowNtdF9H5AlchyntId4Pp
YUrjHek/shYodIKoy5+MuCbL9hTWnAV59DUJ6nreva1C9qewPcEtwelyw053SZgg8bWtRkOX4QUF
qqLqkX1lwpDWz/WBuQPuWhOa7FBMZY3U6fdm83VHNf0+99Av078JpRYJu5j+5A6z2EZDEq41YmKL
C8UgiKFT5+UliRWRfEKVRwAHPb7gFCp2jGyBpeYBQ2RbsK9Ap8FWrbYd9VLBqxRUjdKSOqTmLyvI
BwBMQFZCb/gNGmiZNbzfNU6WM8TV2z+P9ad7RtssIR9cV7ImL7Hcp3V2FrilH+odMwRaiqEj42Hb
tYOTq9DRI0fqBq4gllc3rxn7KLcggMMl2076PlamWXmSreE/+2/l+cQzvCL2gE5VMrgEw8bBQUL3
DIuUw8HbZ71S/ASUsuvfO/EspWNleY5LnyOsz9Ic6x0dcn/veIVHOFMZIz7MIpSfHoD9PeIuphIU
TchKpjylSTqqYcFFTQZuFSD/v+54PhUqT6QDUAl5VPnWqQM5x832nCzTNKI++EelDNsPxC0d2ugQ
m0+VaQjtnzr6eytMhkMoi2b2tDx2k8A9sq5mnVo0XYAvNm7oQ9cMtXjG9/BMsjeCofHd+AJPCVRH
s77B+w7Q1N7vgnRqTteEwAle3LfPqnL7ub9uCf4HS6M1VAvWYfaP4rt6g7krMjMgMb9LBNwCRSH9
1ThKrm9k3hpF6fbzR/FwU+PyCz+/oWIGo3u0E07K6iNr/8WjAiANVZMOa/cDnvs50WOdzsy2XINI
JSVnnonznnI7irrTVioaQkesUdlZODz1Mo0IILn2h46q7mMxlMVsD5LS/XgKaQ0i9eBQ3O3EMMSR
nr4mhSst/Vgb3Qd4sG9XtK30HNdSGz/UKnAcXtrYroF85qTuQmUKEXM6nvKSyeURAw9kguInevYk
pXLhm5AAe93mHXfwp43yrrw30krBy/+GGN41k5uqftUjbDJ33uHduKP0UCh0JqaZAR4qG4oVXify
5mFxDGizX5UtciyWQa3WeM5Tid+m06baUNeGGt+YvWiJEi5QDU8uWCkjyJ38CCQCtPbsN6Jk4sVZ
ogzDcQ4/z21MuESrjI6rZnBxZX2BPwsEHlnPzlKUj+ExWgyqmYuQR0ec2MifDIGLzc2irzKPb1X+
BXaVXOGb1mGXk4EVxUcXK0e8RVFlSNacTWP0GqkqNHQnVOpAAQ/2c64fFB1WusThf2UHq0PkQ8bI
ErmRfxTmlZKv7diwDzio3StaE8PUPPVXLxL5zjowUVmAY01uB5vyoGjohMjl9mleephKM0ovq+vg
NeixdnWBtba4xPXhFKJhA0LE4LZu7t2SQp+uquz8bNRHqG29ss7622t5TnXEI7eIGojWxZ9mzh01
iG2kq7s7gL03qKLcurPFInQ2IHgx1pVUUpgGbBKs90GgkdXdoBAbM/vniCUljD0+79HL2uLggVkf
5Go1WcYEkEceidp5XiwVcT90ZIqkolHDCGZt2WaScqTA7vVTNpvWl+2LO5PWVUBi+Wd152wcQwMw
hDCIZhjfXVl7kpcfN3x5bmGMFt2gBihcBgyUrC/tevaeJtrTnIfBG0Ho/lghllS0fKwrmlL+SK6b
jEk6wy2nlnauiujExCJB3d8A4SpDBus9vQdkNBZHt3vMzYTyHdCrgLhoVJPxx5bV3ButNk7+LCCd
YrfAeBOIlO2aDPeH5sAfdJOTWNpYheNlwiTUHBb7QjVxWcAK3Db8MlDD6gFnteuaFHR/RCwlc502
mPvWe3EYSvrxJFj2kHyPAO6E4ROAIa0GfFGHCb3WZKnHde/ld5J820FDssE+PKDUWjtDYqzI3IrM
uvq1kktq0MifreyZiz51FjKxJeuNQtxZZQub67lVQ4aLBSqFpQkzN2dbUXweJvd73GcZbrRraHqB
dzqQed5QHn/61CgHeqAt45ulyIddoErE6dBrv4WLHNxTWniO/fcECChZ5kEHmo9aD0nO/phU2gOB
l70rdwAYlszxQbYGZkUp0X7lgesiSvedxjdsmnOlXHeOhHmqJAQ2IuasQdOOCTW2PyJo7OBvb//u
as9Z5jf00tauAV5JvBO7LGHradGcUgqcPBNCn6vUJFv0C7Yt+/L9glxvLzxRxmniX3/osvHsEjnC
GNop3G5Upk+3x3GzdYbc53HKSvJJrdv2BaNhkGWVRLnlu7tYFAFA5vhf6C6L6309nRqbsmgV72FN
7JqGF/tQXrdrTpPWre1DQaXddfEQ7RHaJkhQ5GVtxT9ZijqdCQ12JucjT2DmLjwqbJVRV6QID30C
ziNWgJoMKIctSe/C3wtCArhL+ArdwB3ARhXSTHE3IDmrz37j9ihjAfPUFPC2dvtzKhDhZx8oNkPs
7rSA5pO6NXmas7OBjH5qS8awWHenPwIIOz8F9otmHk5Qcd8sLbLrDkYnswhrGhI8/ImZRTO+345J
Gr4hNZSjw5Jq78nID9gSfs3z7cSRWDoFH8kC6gvkK+54Fe10qkPDwKMNF3oOYXhro8Oi23Q3djb2
ORDbydxWNaD2YSX4220eGJNxO96grRlKZgzWClapuCct7L6We1J/HX4poiYc+JWC6aB9ko10q4Dv
eTUdSYf2bdncdHgJ7gfilDzHu83IXZmPEPDEKOaNsqx9Ah5gZxTpPRQRcvkkZ7iUeXRbCzzgoeed
dG4WamOg2DCu+jdeEjf9LYfeaB6xjGGEG4b0RKg0Q2etYClxD2HdNrZf9/SkDoE6CFLmaIrtVCeY
RX0ZVhrYRheVXPENFfQqQjzOk8Gy74c4JUnhAtMBoiWBOJrG0oxQFDCy2yP4swqXY5MnNK4bIagE
udpar+XkhJz5sqy5vEb9ly48gm+y9pbpzqa88tkRdebVERWc9EVHDDknFNEBNOu3NjliOhVh/Dri
O17/RAwrO+Ixave0eOTiHeqt5GqOTK4M/r4ozZlmMaJzLFQfs7M/zDaojH6+trmzBNs4dmWWyOK0
MknXQFxyu+5lRvuDZWK+VsN2EySQOr5jP838fADsAeGh0GMstj2YotaYHkzaaM/Sv4K9LyQz395c
8GdVgqx9P24AGU/4vXI4NSzmSw+2VwaYP6XsiOSmVaW62ZWoJqiHQVEexK5noxNGuDziowfh2m7u
Ut3F/KFihdiNV4swIFI/IrDJ/+eB6BZseSdD1ZHjeSiCNC+W+7Jyvv9QXJ/qKtAmVxrYHLdoJWJH
w8wxdERor8Nu2CR0izKZfQw2Z8Gv1EqdYu1zas3LxOFN2zQxTtSy8oZoz1FZViuEUuuhSEYIy1gr
bMGZg19gqOumU/SyDWbIAMOPs/jeVOOn8CYyEpsELdqK1isPE6XBw0sw00fSEHnLb67+OPhlvsKl
1TQzbKhHI+9aUraRneLkKH5UjRpnTTbw3bP0JaW4aDQ2j25gHL4hnZ21UC5s3NYbj8KcF4gYfpbn
jjVwKkHswXi8TQ3LqzDH5n07KupMtzu5u54iyddSBWDWVb+PiOhwdL66O/hjzWQhFo2VHHViRAkG
oqtTsUBq59AFEvIOcL1jnCMyIdL+52/qrPCuAKbjpfGNg9Rhys2Hke0eohUDNEf747F6nlUEpPnz
W5Erug0b1jrvRF8+jixG4kL61NN7bm+t8F5fTymbxgR+cA4xPaGM8H9qHLahUqSCFRDt4i4wMLh0
I5fQF3kz7jlh03GD3F8Ra4j5u7DtseQ6jk6gRLSqw/QgrJDtNrr+XqTq6Zvo2iiP8W1dSIb07ABk
M8idKfbIKhfYO0xs6ucMGob34xCm4eLp0GPyJ7fiTIMs1VahP1arTD1v2VBZh+qvQYjBh4YiHWFI
agp/qClxlxz6T5QJ72BPHaWHXVAl6MdkkOKrXroTPpU0kxNvg2wHnOox0uUJY5rhrIuaoHUYJq+h
6+PEecYUTpt+mAOuOOyYa7bnGftyxtO4VqbCLYccHGxwCd12FY7nuwvuPDMtTOup8b44dNqqqaoQ
JdP4Iy8ofuz5J4jNxu7tiY6g/v88UwDiFn9li8dWwsj7e6ZxRRba4ZeQz82OpiT+uuH759yf4Mva
N2HQMHCkrpTndRxZdEscfIom1w41AJur4WcRl277ZcyB54LpZC40Glm12GJh5LQkvXGO/IwJKZ3D
Ut8MKkiS4XMM6nQK8z82xVnE9cLHDHTfwYuc6LPMpLi2Tcqa1V804CkOx79v40fIud00cZx7HRqt
sZrW2TBtGQB5Ngl/Wl+EBr+//aLk54ox7kI7g7ZN71U0WK8aexWtRuFdXcUG5bQVxTzCm7fYIp9y
0eBCuDsSKk++tLumLFpW2AmV3yhi5t7v9oaHjMPidH+vx7n56v/0SQAfWyFuCWjZldNwzVO8BdE+
I1x+TGNbY9bn0ipKK9BU4jA9WY5ggWWHqvmxhfgHXHtDhVNrNgYwu5D23u2CS1qKwVYmNEUArExc
9jt1oa1IettKpWzJ4pcQh6dlMZlKTIQWPUdjoqIFuO0iq8DOnsgnOQeU4MnCcwrB3rCkyoeBXxRC
HMQo7EU9K/KcGQyg+Taq54eg0E66v6X7Y3bbDJt6OMDVSQ7R+j66Ge4QDfkMVwdOBHw/IWfvMWKs
EISvRlRRB9ROvxzIQPfDIaO22NndRsGJHM6mhdZUi8LHn4beQnR62Tn6jHtwMfQTd+dVX/dGB+jM
fS4o99/PC+tzFZhgBgUmrtLOVZRB5SOOSWnhBUrbLEwzkWLNrKnbz24jRqiFh0NNyj9raYVT16qy
4EGPeI7WsFb7xIDitjOACdQygMM6ZG94lVphq2B1O1xvCZ+L36HqDz5uzkNJCCcsXz7pm4fmYxtt
m62BdcK1vvTGV59WLvdt0/XjqNXSpdzaMYxLC2w2VeeA7ua1JtCn9tPL5CtJwsUjV5p1f9+GPCaN
Hvmo8ndUKt0jy9IXxJb1EdOy25nXZx1Mdz5g1MR0G64okeKtJwv7e0+LAmtnVFQHuDx9fmYIaXtx
A3hhT3ut8O7+uCFAkRFl6pxIRJjwBH9ZEIAdBAD+klry7s0E/CzeVfID4pkCLbObIYtB6eAnQk6U
ZsXyLY55ttIEVi6ZRda41S3zW3LQpsZhUClN2ESfWv+Q5U32gKYtR6dnGgZvCnqTRQ6cdvBCHZh1
lMyWy9s0TZFHfSqeGRYu1U3qaFbTGmguq37VY8G6bc6SWXWmUYdTjP2D61WqLGxBulGYLFg4Y7Bb
87M1F5/sFHYO+BdefveZaZw/xHGgly5WJM0exBYIkUQ9liYj86vWtpOzrI6gJ0mzitWmog2X6UPA
HOGn70+rFqVFQaVpzIZ/y43uk1rnI2j/3CLjUsJ1weZNuNQr+gzRLXPcuufWP5eeaek+CUyARS4G
rw8qJeE/c+by8uvFyfLC7CMdYQHJNtFJNSZFO9hUF+fwDnhSnldyw9EnL6PZC14GLHmqQpdS9uPG
/tzbWFIA7x8Lm010XXv+Wh71eCWyK3IXEFlmRQ04Qb2zHGf0G9k44HhalTOVgX6m1A3NpDdZ9F0l
GEvFug/kYcLNb6x7sw1lvV+/o1fqrdrtZ/TXQNhsATLTKGOZ+HzX2a0z1n3BNbPQKjOoosMp4wI4
Oui3bbvR7HwCVjTRTV46ZqIG+AOAG5FPviKSyOhxMij0z/RE14OMOW2NKr4Zai4Swp62FK69LzS4
5uBBHie4XX8D3ine3QNowdAnhNiACmw5qcTn4Svc8ta/ytHsvTI/oVCrO6gEh9h6XbMzr8d5AYB0
Vky05s4YQylcMx+bJZnCqRX7u8UX8r7Y9nBAQILhrtdHO8/O1/iS5x7eIRCAuQWFLI0nZppjyXlO
8i+3dfyRxIMqvFfaIfIQcTzHnDOPdLbNAEPY/4EpK+1EsMHErDoMdGv5MZJxQo6u3VvqTsMZ6lL7
hsDeM5rNz7CWaKDvciH+oRMdTKdQLP+7o+dBvNUB3r+nhVhc/BT2hjUCEpF2mK7HM0/MQAzCRDwb
D3oWeVT76hC1Muk13V9E0CAMuf8fk2XDX9hvCL55l+To4DYhoSqiEf1qY76SQR7p+PwLMYiTjRwo
juhz/4zs7TCWim6v/ox8lP1p3qkeoO7zsI6JwACJPU/iJP1Wwc/iGL5plRUapYdkzK/pgXdJqIyK
lNHerzJnlrVhFc0zlKpqbYavCxi9dtSp+X9xXifaQzuwL/El9BH1MxksWr2hBQlP0Xao8JHbB0cq
Za2dvKW2xzZXvQn1CKPg+9tsSBUHZc6XVEsAHEBNO/XBmW5rQOzHyMClU66q4t/z3GHEd1aLCPFW
6wDCY7oWyFOD4YCxkV2yCWbl56PfM1pTp3j1rvkG24yiQPbfgc++holpgi4mYKhgryu2V4VXd2aH
QXWOrpyPPDDqgL1YIT5FT+8eXH6KBVmkEacUxoPZ0ldfXKGzpZKLUSm/zYacHviPxIKLF6aSxQ+v
NOVtuKYiuCDaA9g3rS/4vtMNvfxVBaVXZbXVM7ZeOh/o2kA8lAuPcaVxAaAuYvxJUMgb15nwwe5F
E6rxKa/6fCqXKfV8xG1dabQOIpws+agGJXZ7o92DFIkgCzzv7ggd0FpLyzFW0vA3Y7GVyg0UZP7i
6qgr1jApgLBbt8UXfZBXClDw8RVxE/5nj5rOy0HpudAmEF39ofHoCYrrKTjpEIS0JmBC0ePHewZ5
oTFZniEIdTvgJZx7HPEm3y/sqqtXdur5kIym/bcngma5mW+rso3aT9TcMyqNn2hexY3tNHP53rye
ao50QeJ5FdyMErfvMQDl89caSFO6E/Arz6H+JgMW7la6jDbqB1H3VTlYoalaTDcFXlE6Qm5CdA00
LxquZyv9B1HOGBQ0fpcaceO+3xDDwtCUL+TZBkzIxlIvsArrD7aI5KmmnnV95he1stiNUoBjnj0K
h2/OjTulUBeTVCgNA81WplEFViHVaVZ33X3KorhA2+8AEabt/AO8L8uykUn0yUQaGO2olZAQDSBf
lVx0KWbtUQ9tcwx0b2wH39BGtlfvpb2Fa0HreztDalouIXxiFovFHIjl98mt0igORh77ZS6ZNJDq
QKiSP18kAljMnl3F1yC5X7lKcoIsndn8+zZjGoeTrRWcDCR1C4azzWPLqBPWgcJsekSTc2qAKxOa
TJPgWEHoalYgPpD9n+fJXYWN5qJ3o5D/RkSWyx3qWsconR7SVBNCZH4tFuWHJ+BjhLduhl+7RGME
QkTqW3YIRsYsRuV50Wb7gnhooDKvWP3bubsRLoJAdkHZVAuLGb9f3tnM4JxEtcjFWgbhRu4pCybd
utbpK2aMQWoq0ZUc3CT1b1bXRG3K+js3XVRkbs7Sc5lhZXFLO+/52vkOrOg+otSt64Ci/dZtV/8V
Skob5BYXWodwdZSTsGmZH5IWM8Ih6yyrKTe1GH1xicESR30P8p1sMx8muCsMAnpDSwihX0MBgwOK
taaX6wUJcFILmhI+AVlmt0szoJCR4cWHg0oql/tTakqrqC6/Apnko1svQaKi2+mbiJdbULbrOY4z
f70Z5s1fDpKBM0elqD1dZCgQJ7f52Q1nGZXckr9SIC3ojjZvgz8XQHcBozy5fXjNGkzWBwCjPq+D
PkPpJBMG8qWe7fdFMlHhOdJDZ/ltyw8uVS1libffMFEDwTz41H7b1jRtZJfDyFpI1V3406/96EmR
oRE77EZqnQ9WdIY6DvlP4uh3/y+MCHrZLBblqZorGtKftPxSlXY31cnTADBy3txILGoar8cdah8C
KSOXMnh/BT6GQISZtWt7zWo5AzjgPksihUWopsMl9EkSr1+/nDFlKEAZ49bOPjlofkr8UUqeqiDe
hC68VlKBc6TpTLKzb0wiyPOFSS9PjdMbxOPQkgNB1+oV0VGGSSrkdPX3pB4Q7yjCO+j/k3XP33Br
wX/6GHqkAddsv5t0CoM5+5Y9gLqtaE9A9bPqaPTAB18jDBAkum4lTF3bSJyIJ1WulRwcl3OtPBcE
AybNWwUyiG4gcKkSIP1vzBf9IiknLBpLbT9Gamv6q8mhNoYxbX9yq8k3eVW2M1IzJWHIZP5ZlT5D
diDUBb7hZQccJSZyANvDdv4YhPmQoPK/7PE09Q5vZ5H5TzdOriztVnSo8It74X8siuixSiiR9Rqs
OV9g2sADQ5TDMqwt1aMcLdy2F623qFmLhL7TQdQ8KwklU9e+b8w5i3p28DcfaeJG9x27jDkClfJ6
2v68v8WXMnwajZIns1ChBKUQvLAyoN9s5Slw17iJd1YdGvFqiq7okLC4yWpHq1CP3ePPXJzWW3xq
7uyuPDH/7J6cyNWT8sxoy5WiXJDws6/1OR1Df6SOkYBQYXcQldV4BzSWRZEa0EFUcljW2HklLbQm
5pKuQZWxh0GqRqnWHhx1d4gkCkG9AARVGHtRK4OwUMP06KV/6X35AHmsvEsntA962w6uxAMhng7K
iiQxB4xbwNll17beScbFzObF2WM9kUIl6FXFhE2uK6o7Ssd4RxH3IBK/xQ85QIZ8stcL+NGcUvb2
cFHYQRZQlvhmWFtF5ne6ZFxPnDpERVtzA9fRs8AkILY29lJVrYOBpigTlZE0DjYZPZ5CXCfApixI
opO8nwZhiCoI17es7MW7pBRqriFJP7+blvQ89tPWqAwGlaQsSPORDfmUxmebugsaY5fnwR0Ft8yW
0IMu8rmgSq/CtM+VS0Yr17gI8b6hFePoSSwIr1DtjPT+E4Y0TQakcXaDecAsg+2bFNWB3nY0rZFo
QZ9d3dS5h8qZQh5LCMYkoUISuqior8ibOlgvJt2iWYYM7/EQqQMXhItLVnlq1b2wH7LEliNeMtNO
ey0poZgmbfqahi08QXJqnYSiF+3T5VCkCCLYGcR1URXHTxmcvb+4VwyFhIXyxz597modreuxawSw
FmRK/BouWAWf67H24HlI7Vyu5lJ199NEP2Zx4TnLJwPzd7eR5po0vbq9lIYDU2mWWvAj9Ejo4fHj
KQkzdVuiNAo7VvR0x/wPk9J1vhh/fcRwPNQkcr+6WqD0M5qQ0vGJF4PdwTri1OHEzyGO8pbTkGFU
K2v0CYNobWFeVkQcfdyViJcqhYEn0eGQj6CtujrT3mnFiWRR66xsXostkz9Zy4JOwM41YWe49mDJ
xwqeZhng0ttJrWk9qr2mlOTt7Y7E6haDZ5WL+6QOuN/XCszu3Z4ek/ud846+SsVbrSew4AS9CcYk
qimeAWf2m2CpZDubRvQUELhRlMvOAg6gYa2tx9gKTh1usQrBv2TymJV3yqyGh3olG04TV1fR3VL1
+o929gw2NbAiN/9bJ43MLdyBSGZALnJCnWss2jL4vOuvDR7QmVzAkLOBl/do0cNmrjBKZ1nsArUu
BWVcZM3l7/KA98L81g6nls9gJ/4hBCO4HR5BI/t9nIhWt7i+axrM+DYEOvgewaExd79Xw1+62gTa
5SfJ6fQmqcrrUnBgZJfOw30AfyKhZ8pnI8sGRDfUHkg5yJp+FvbP0y+q6X+5vQFzNVccdHvCihQt
eJc3pBefUsYxL5YXkynhHvSX7INlOyI0KA4QG+UGVfxKBYaKZeRbkc7EGIDEQqlbFXVSHKcxcNQe
qpcLXFXVXYxXP2oH2A3xj/RwzBVFvXqXqbC/M5y0xO4uu2tCwsVg8UCIDLzuvZYztaJv6zvo9vJd
+n8yQcY5x5iAQTw9fXad2L0/ppJGL3E3VlYXkeLhpIWbR3RAs8tH3sELazoPhvm7sHKWLpkmwP6X
6uhDDkVc1DJyNlNOfaGxXraiy/ASt5HRS4fTF9uoibFKSYIsgxU3UcZ/tLp97tFvXT8RCNXJWkPk
thdYG2BSi0OsnsUjImkMwuV3KEYtR4V6ZkmxDHM8tjreAkAXXjROuvTkUuewTjO2/Rd2rSAr/Ry3
9zpoJXcSSOXFmWRAU3zihNf1mH3TJu7rLSWNUZzgRzlNEDZKcsdYIPtcDGY933sH9bivK7oyYCYt
wgq0E9ewTYxenjr1wydNH3qtd4rG8/o0StUQc7kLzg0mjEUsOmpzPoXGVFodHGEPV4zeDJqz/CxD
VMDGJN+iFhjMSGtqdSUaTMjzy4blpYoid+y+Wvb3Go9K9kTWbC2FqM5MlHuHMI/6UrzXQ3UaLwIv
coIx/zhk4QHAVna2vMJJFBX8bjFsyw+brgyst6StjgWnXIR+BC373NysejmjNinJiyLByCWts8Ng
AVz1XASXhvkJGaNzrWjPfKvVX7Rsg2ryrbZWFFAIGyvtq96CYnQwKK3xSQNUoCQBxirl6I+FqBzN
8vMzkeMDZ9rpZbdR8NobvjxR7aJEWufpZBG0gcJtY3VWhx42HjEOHJbvJzn24jBwrn1qKbMDfcBL
hITmBiPa5WTGC9cimK+bpvPs+/Mxy2jln4KGbEWMhOyeROt5D8UTQDlZ1rqyXD3rIYgHrmzoYn/g
tqD6Owk7h5f70Cwioy5w75YSQbi3aP1y+UYwCy/X45uhwCogaho2PBR8L3jFm5cDYX2SUMEOpVfU
SM2Q49DhL7WwPNwosjfS3v81rp4O15yWvcLKputvUfY/2NpF0ei3Ml2RiM/IjCqVxiK/nr/h6fXL
LxPuaUb2CE/jI4RatjUuGzhKrKllr9I+CXUPIoGfZCpHaWbny4G3PoKVo95hzTqDiOLVr7psSfKH
GTjGfrZmOa0T9OjxOmfaBxdqyomCw9mUdPV19n6cUmt/fH1YJtQwaykjUfndfWkZ2ulf/g4gGrX1
+cQKuaa3Aqg2Ff8k2G+Fev2AeMHI0sPtABSrwVUDQp6Qv/fzSYYfGgW4rALawde6eanxS8q1alLB
ingumo861A4WMVPisDTW/r4Fu2/PCUJ1ineqcxB7FS8XQddIcBwfsiZcXaEkpCBXQ0Q+7gMozcr4
OWvUVMWsa2qGHin6R9PDejnMiD6sLFVDXlPK2nWjAglMLVrS7OMo1rxICMqt20DVUc4Bi7yvPjHh
/B88H+9MRY2Uv74i4KzKHx1v/JcnELoK+UKrbyV/bjdOXwXGVCR53LKJeLG8yUPyXhw+eizyKpqU
3jXM2gpc4g7MYb4tU61Jnfp5/UN00Z23m6DKO9zsDyiEk54xrfVk7ZcrkqWkavBSSxUkSaeeOtKy
ehSxT6GyGWw2sDPS4tcjQJb3k+ADXArUCoW3GXlUxflbI+SnXj5k17oNNpestHCsYJuCBNgkhIbe
OzCSwN9CkI02R1KdhBfRB8RvXO7my7E7PFn3Q1+JYJ+p+nMDqbHXpRjTSCHqtfd5bFAUQQbv1US5
fOEmK0ae5pupwtDWCSQSNHcein7mFNKWugkxlsA7nG7OToQWNqYKxIQOY1ppwwUL9/N1zSNwIf0D
6iTqZZmxpFBFChuO9t9z+Cd+c2KMQ+PTvOQOS6r0IVFE7ytit7rxfxZNqESFJnvltlLbb/O06DUn
XcDjavh7CHOe6U3xByjwxASSLkDS0ylpAgiS0QQ7IEM50Yt1x81hvCSrknRa16z8OHsq6BBRGfqV
sdoZEm2zHG7kKnTQbYqfw//51/mBPhPNpRI4CCxsS9Q2UDbd79scjgebbEeJx5hMceDV4oYMg0rx
FtfH1o3X7IZXdRt487bitmSy9RKmO+pHU4P670PFJzmdzHJfVGKjhR9wZ3C8ibqgPbmape4X0WIV
c2HWbOd91OA8tIxFQm2vn84wXEh08BJ/e4VWQtgbwmp3izWWwB0k6eBbRkYFb2ofhqlYMqrEZDUP
IAV+lcb9KCL6txlO4L5syhUkUhf69ktpT33Lcn3ZWFuIPJ1wVen1MEIafIS6s4HYKDkHxZjn2V9S
Ap9X1fsnNcWbB9qNBNZmAm3FiD8rrA5dRW4PUnmL47fCDXrvXWltsREtASRCwzIhDs5V3x18fe24
IkwYEq1u5b6mYs4vthBPP38RPwO+4W4Ang//rHKsy0Wnx6JA2ZKtX9FzADWn1bT8KxbdLoxLossx
JdFgSCxmXsQ8xgtqN/IicvfPUTlOdaIhKDjuKYrZYnKKQPcYqVkUwDp0qTnHE0qIL+ty8eZCzGcG
SAZcJOEUAnzfMrR9QZsxKN6jbADoRXFgwv6gL3nMwIYB3yi2emuYdi9e6gNPHkzZbplDgrrrcm+E
rh5y2wIiJrj9r3p8oZB7FjKYR1IBQtRy7DQQG/8d/QwIhwWvp4S8yOaarMnnHazdOsSrvGHghmho
GjVjQ8jzGc990Vbn99u5U8w1cX15HvYAEeGb26QnEFJ1XTq/h7TH+HRFs6jVbkodDTK9e4Jaz7jr
2wmrGV60GwXwSOJDpKvsvKkG6tOUWLV9rC251vSEffdySZd2IkVqQm2WjdAxMzrvA9Vr4ausJHsu
US3jARYFwuMSyMipcN+7UCVxz9Q6eYLn5ZaCau1BudosIaGVQ9GWAUh0aOEDAq68Rqqqn35GmI2s
uogamF3xU1Mjp3A2PCyUlRqwj90Tk/LP1KZyc50JCY8mnmNhefJ5md+hdKCovohZ78rGtw/Fqxpv
UPv8HV9uJfa24L8U+Xpw+Wl0w7Id+gzWNOQ5lOZMGqP1d28O4cXv+/oW2q2hLUbIYwyfl8hYAF20
jCjmmwyQ4TF+LBf9flLyvVikbkzGd5tUEX8221sJWboZxwGBg8SWxqTdIKXN2CQUV+4QnJNnshgj
KgG2tNJBBHDrIT0TT4Oh+JOSb/e6yYDHEme4At8rXRmCuPR+rSoEEmmgBLPbRoWk/aM2ugyZtnEc
jKCJj7m2y9yalEI0tEX28G8UgnvIjk5s8aaAP8hn++9J3j30req6aUnYFyHJKIb9Ueekp0JMeyb9
vNPjOtMP10HF2ny7NEfueqdW63U+1rcOBYVBRt2w2CoEb4UT0Z/zxqJuvLhjmQ8y7+3GYil+tTKr
VU2GpG9w00rZIkNFyJWLfUnznGHYLFhGTot+tgMnNG05x8jksdnCIYztM8KJNHM4QZq5Uay4A8sB
cHkJCvz/x2yuofYd0vmvgH5TTJ8fTfPjL2UhUY7c7deWtKG0AxFfu3M7hUmPRZfnxr0i95FW/Y9b
6SC4+FM8Z4S+FmcXOFIjMZMLbdZBlyMzeDRCMGNiPsCz9vryKvjKnJCajc/aBzKj5SK0rKSQu6YC
jwx5z64ECLbabggsJsxlT/gF4CtBphG5ayTeR/A/8to4d2+HyAn1ZO9OrJnHaNmn0a8AliShnpEw
DEywyTiR5qoqBZzdehMeDzscswd7BPCfahVzdOPsiuN7k6dCuBr1FwH/hjQ51cfKqm61b/EoWqFY
e95b6V2rHxdOvFWiW60MdJWaBSiA79I9Qnfxfbt+thPvdenyt01XWgrVCHg9uwgNwBR+LnILsHlF
OZiM92OvBjcGY2feyhhqCoB2eL6OmuL5wGU+nxWwlw7e4sptj+x1w98gXN/xSvycXpWqFQ6GndNK
K6zmj0/qXdfmLyut8vdJJ+0VjJaPE/hlMhkAea60EZYR+UHqRN9gBkADMlK1YvQ0h3IUXFJxAdEQ
1dEr6dhhaD5K/+a51rLx3kAc5pEgp2nTRPo5wV1iRcwfV/FAul/XUNew11Xy6Xf5uebTek9GkU0O
3pQam7rvAxasY3zDFarTZxSu5I259l9m8snf7B1tjViqXH/9GSy+ovMbsUt7LdzDK+4RUudVKJVa
8HODIiveF+A335+wL1V2vzkCCEmjzbAW+htt1rAJCXfeTKMZiICah/ud+h9RZbZAhx+Nv5p//dNE
Vd4XNeyxcpoVxd+pfjwvo2nkWKEs4FSYv2czdbw1gfr4UPqnyGqFexhrJaK8MBZrsYSerhJeopxz
BnDuKFcUD7ed2Omj2kBL+5kN/YDqLy2z3EiI3xwt5i6UqJb12emtK/l0+f25hna3my9har9VBvs5
3B7Ms9LROzrmCeRI7kCQchqmxyOYyItPnBPAAHPgvIiZvDIy9buS1LBESeuxRwiJpFDXzAEWB/hx
cH2z5lG7J0nknZeb2StyseRULxUD9M5tuzrZZw4YcBacOsqMUILxUnnDwdViQUNTgHmkTxvAEToE
3ux3oft5C68b4yvcqfL/viaQijaMyEtmvZr71alk220coEhkeJuFwzEnxjRsHm2g7BeDUBJKRJ+V
Kt4UeePClXGRPQy0gB+W1Itk4ykOLCTtWMtVspOfQt6jMxui4ekTNDWlbn5rukHlZF9tNdirNRl8
wRyatof2PpGQRAz5/wqX0y53TSkCc1v7AQ9Oy/+euhk9ZPDmxqTec95VwTbKla6hIYDI5+PO4gca
zlqoEl89JqZjtl0AYwU0QF2cZukHiRnh982SYi7vGBkoTbauF7V3f9zgy54bKmX3icwlx2q6bR1u
nyNwVvnP8YHkJiygKcTRD3YtnDvJ7YceOp95MArcM6DSxrBoVBDenRPeRQGoPUkwPEHPick77rit
esnC7q5HEv83pJa/YE8MRrWOrK3TEhCkardp3F+BGqUkqd6qZxT8amUc2JRInMswwYIoz6+wD8a9
oZ2vTvFDJui8JfHP4I/u7ap3MPuIYunGrMk6AbvwQSfbL7UcW1j9hvD4cgOnSRJtU/fu+qKxi+bp
tjAIdA2qSwN+Pz92w/9y8z9UHziUjCkUc16PY55vybcvvYddaWA+pxnZwGcoe7zZ1nG8PJJZ5OOr
fCBK/ndg3OPSx0p+VK0EyKDsigKpBUpRXo8wq3fyokMo/vsN0LfnPIts87Xo/YVzMaDV3ttQn22s
61isKdrkyiKUDbCBwkUHS6J5SIr3Ll9VVBA4oGM+OVnrp2QxyovIKnjG2W/5vDgpYq98KLT0jID7
TieYk7eW1f4uIXF/dDz40OuLgZurbwL2dY5R2V4IqnnlqWZhb3x1oDk9hwFUynq7Y9TpnRuyJpLV
Qcf/QXDBX7vrdEJPJknaEzzJrXCGrOqkFDSQhLS15mNXtc7WA1pDdNikHlAcDu38k92HXrjE0hfN
943+DA1dQk5vp2lg91SkvSzKy/NZuLWnGUhhOZ6tMGikAOs12oqlyk/4qcyC98HDA7J3/EPIS1ew
dmZIcvebi84ceZq8Vo0cLHM8ffHYdCxNZtj+j2kpyD0+EUl9NZA2SDgey5T2+YkEQWorPQEhdwYY
zEmu5OpKt+5rMpUhm/Hq45p2T1/v/NjXWu1k3aEBNKuQv4TgkjD5XY6TkQz5VAypfjSHQ0THfFIM
RmhVa/IN8CoaxxakUus9XQqJUppdeJkaA7nCwC/+V+cdxKuo2buP09wqBJHM0P8EY8htPI4RdZly
nk0gI1U95LzN+/Qu9RHCumLgZpzbO+PH0zvyBZ1R3nXd3+yjMPcRhaA3BHK825PDrdTVZXRBEeA+
rqtJrK5dlBIEjAcGTI+Hpxv7CR/FI5hPsKN2PmSBvq30OPBtydRsF9uJVzE1pQfdf1c/vkrsSPjG
LUYN0EFP4nYW3b/t85mRY0rWkgwXoxctoRf1vEpltfYmAIp+b34XQ1suCR3swkqZzSU4r+Chcgi6
7N4jLu/f0M1EitXkJtzyt9lXJTha8PTj8JlHYtp7cKTF8BKGywtjYqqcho8S7rZu3lVWVaihZeXZ
36MmgVlF4qifJ0SWEfh+BHrb4cPZKp5DL2Ya5mEnm0vuJnkXNbmH9lVvs6PWXNaAK3lbEMxLVFLH
IcqFtggVOLQuXv/V+gt4L4smk9lm/pSyLmIAb1LBOCjxsN4q/zwQacqvbwOWG6o8pM2w2SdY00EL
2ueiKHruS5SPE29jrCR/dYWvUZ5P9Z31fbMRWyFqMsIULMChhSsNg4FIOAABdyb2KwMS/gBv7AOL
g878HnDWn+1ZdVowPkz725ExI+Btycrvrfbj2mFljEJv2sfnAhW1Bz5scMU/Le4PvOZkcqVrYsyR
kmH8zUq1QYOCJHS6SVIMl58l+I/cLlVxkEgNIhfcagACgWvNVDMsBbnsW7J38eZbwdghPCqUJYUr
0qyYQoaMMdt10ruaCfA+a8LVAR88DyXquUzufM8aGLdlj0pOqL+jX9rUei/jTVso9aktHOCMyXEW
NQiv1DEpcXOxKeiNizxh0P9foeGr40dvqdGf9/BfqaQLZLvKd66HlGohnStqs4MW0RA2/VBW3QhH
UQmeU0en1p1hOuQl9lRo7ucaXWGGu8eIF64SRUDwedRaw0m9HIMsRP6+OpT9z8XUZqcxv3je4fZn
Dpk/fcFJyG4uQM1Sf9L3V0pddlRiDzxTRuLJmh3JtKt/YU0tasqphhX7V4L9awgpow8PstJlnySa
ARNg2pvtfwEpPhMOsUNiwkIwZbYzYRqAt6Ax19mpj+KYJJvBH4ZV3cY+0MfNufwczI0R6MmK/tKw
XF7w0OdGuhWUwyx4Jjjb/mRMgzCOxl5DLTvtBn5tE/T7gzGdpgXD5gH+5oEiv1+1AbZcV4qIz7je
edQgG+kAjefpBIuUww4WcQW27oK0naK47nkmuW+vo/CVykueLs04npMdqe/nTRwalXtd1O7mOgis
wwQgcL19DRWiyOaOSP/9MAf5daKYdmHDEXLptlAGGt0B6XD1MkSprWC/A6lRtVEdHeLnmC9fJo/q
rfaRDphNFfGPHp3JfNUXzXbEED60+iJ8o3DuLsBWRYHF4Gy10FnXTp8En/m0PfNaxN1VyrtnlAZ2
oTWfmaDn8bwxrsFpozh5ZXNzfw3lhA4RY+F0taeMJZ21LR4zmT4Qey2Pq5RA7Ez9CqG5g1mxeINn
Vkhu/If9hLz5q7Q/eXYkyZsPFTSpzYH2z8kGp08R30UjyqfmC/i3XQcKCoCAWLi5+SKkoHPIqb48
6xZXhaoqHMleIN8zswosywhRs/JDgfY2fEo0lSWKY+PG0fqC4zIC1zgFZPgD1n5uXnb+WsKJcBe+
9jLQASpu2LD3gEvplAwbPI9jR9JTx0O3JyQ56cE/c8HJ4H1uG15S6mt7zDsUvhaZAt0zryY0Ybwm
ElUFyXRtK/2qdI5Z5mAA2DMQXlWrhSSdFlyHw2TazseTvKBIQw4fnYkBEd1zmqPbNNPb9/5Nrr1E
D6fB4dXYDbCMVP/X1scRjov7mK4OdcB3u05dlo9Y630/523xz2Tzyj/KV2+ZjnPMq7Vke1Y20yGS
1/gpebjaNsLKmgX6B5PLtBsBZltc+I8VRFENBdqJeI01hF5kHoFwrNfpoepBZvTl/d5SPVRxuiAX
ZgzP+o9bGjRvubdaY1TKVZbdMtZk5yznfJP5rtt/r3POJb8SeDi4o9hB+J9gtJsBDP/JsInskr/W
p4SEAxmr/WimunGnUm08r5H5j0bmP5uoUBI1dfGjN7XKIzOvcK0DvN1+vCktDPrRnSyeq/H/g+sr
8hqlko8Rbg1rCzpccrrff9wiXTM3QN4Prc51XPH1KqDMC8AqvC0Qr2QZUqjYb8LaMzDoRHXk08ZI
aQLAnflbUHWukCxXQH8nhTdos72C/C6PoCw430QENiiVtCjNvjG2kUCU5SRKV6F8uarHBVWDLqqK
F6wKCjjILbPPcEpY4s8LarXxEEYoX2HSxb/Mr34N+BIM/amjJ2f1zN6oOdEgRnwLdKJcVUAbxoPC
QM1IcOYbIqRZECeXnWdQ3f6/DPEEps8pLnndrN5CHjthDL4xh2DgaAEvDxWe18vGlXL/5obsjK2z
Y7904bWtAqonC8O8G6GKIX8UtEjOjoaAAGqD8xL+YLzXlzA9yfXG1UCmw4TJAevKAMJQl71MZr1p
68z3TzgJXQsDTsORl8RRSILj7iWQ1w0XswwODevXuttf053sZrmT5WOa3SL/VEOCMxc9xGhbYxuW
O6i51nPka1RwzvJDjRHQKRu4mG8rT+qxFPgg8qCm0bVGpzjIffkmK0WdfE9UjRAhG6jd8vtjjOF4
YvZAocyi+Cipb5odv15hLXB2CHuKaHbYLb1h8WpjP0BF4J9XKfYP6W70Lle1oYFaCjVPMo02oGxG
Sp2F5K3Eo7UmX6WsFe0IIu8BcEzYXy4wZKF0QP5n7UcqRos5TMPQ7T5IPeWgy+vg9hWVNfoPwQet
Db+wBwjGBNrygIG7L3neso0lwxDSpk2brLVNhtBuzTqeVVD2knLOXf7vaW82oMFWZUWxAZnSdM+r
ECsmHjKzy/msjJBszF7HUtlupDLcXmOMADSdxGYtgH8IVvYJ8513bXpeJzRDkn3vPYdRXUNNJAVz
S73FtJQDZryK+UG3CCMFabfeWtGxDcZfpuZ/XXQ75CAx/wNBD/+r9H1oKAyWO/xVjWC9iizV+EEe
gvc/IcJjpx0oumGARx2+PRSj9IJx8hOsXXBZ3HDU2DUPsbhIBfpCk/nfWg29vwzVC5cF48154g2G
elRldSuc+L9tRUzVCljPqHpe/e0lspFXPWxQJDNFK0uvGhkfxndgARu1FktabGW3WPbSU1cM8GPM
x9WS1/W/VGctN3q49AvBWxXLx0ERumQkA2PUn7vr8yk6xOq9MmYaD2IXqi5xrfa+PxXjsabVKGkI
GRmXqkBnmnYJogr3TGTs9kzJb1GsxnrXUkL4iBuBdCFOUxFq5CQpqCBM2D+i2Zm9SA4qqbtB46Yv
+YNjOt69wDUKo+HSofOXltSXFq5pMIIRqQBGTN+P/ZUh7ubD+sEw1YVad0eCSNcAfoF+BifunT/T
UuoI0Pq0YCZmd+9eI+teYqHmp/IauZQnCKPKc21rIHaQBky1fnD7fV3WAM1gorqxgcOFwa0V015M
GJiBCnS5FCZTv/9fiExZHAQ4MuezcYcohBvW9X0fcO1dqjL7Ji4vfWfRCYSv3cVVy2ll3hMhLsGE
gndJ+GMwfDCj2P1jGtJXbbErE2ygD/t1VY68x90aswljTRlCEDo6MS+MhAnYNwijRMpeRw2KNsAS
oEbWvcpUQdLejCmlbHQa7BZ3ydtGWIf70fYD4zOCSIg3YicPKxgeXs+pG+RyoK7dRF+OzYgil97A
YN+9f49E9wTJyFz2hetHaa4MiXKbcU62Oho6AfYT9L1cHIzPVRvCUarfBjJc90kewnvoVI9FX/a2
M44Ok9jQJbQAha66FlAChUnPM58PwDW0iaXGSr77vZpW2z9Fr9MgrZfebMSAnwYHo4uoe7Dbf7Ku
h+r8G1lik4BTKBxZ9kFqEE3kzc1jJZx4VKhLUN9t0UAkgYtMKoumdqIAWCaR9ZS1mdZC59OnOMgt
v/XeGv2+/MqqFVVuzSbk+y2LMt9hWk7G4XDuTRRMeTMGU9vrmYfwCI3folkLLu/hho7rubAf8A6f
yXpjxsn8DyCnt9lCoQr8UBIf2kYd3lFgi3mQINmzl2AxoPEVwSUcIRdMr8rLexycQH/LpabHL2g7
hVHUkaqympXpWnii9iSbPKg2IehTDx62lm9pKjSokGw5XtubMC8kWCDuOPIquAcfcw7AYuEXhpZQ
ZickhyfW+ePcWkSocJl0aLNGwOiSlkFeU4gkVrurg/j5Vt2Dzs0dqG7KSIlZ/pk+/q+gNT/yXod0
OsoLCb/wQUhODUBE9OsUJxaxkGJiJCmAnPjbfOTDTjaIbJUfL4ye8wr2mWc+i6rHmIMGKBB08zit
2Vj0uhDsaXjmvT0Ly6jIMY0vfgH0PG9KJYhasvtdrS+sUULFAHcsBhydyCofV333Ivi7qVXVSqa0
ZkCRttWDkN4yooEDWvmcHJjKZhCvG/SupGpeWemEKzZBeaYtEA96il/9cTKHAvwJO2UFg4yHU98i
IFtiqbwKF6NcFnZcw3YqTvgjHJ1zueGjsVODVtIUYtc0Uw8hhmf39p/iSefuN+DBEaZ/qVJSUVJo
4nLS0pgFyO3KRhK1JuK05DYENtPwH3TSDoqUmO6abs7qaukDTqho7lhP5gBhsGZbP1ohXEM7rUTV
kLl+WAtXuAtuKpt4/OCPWZYEZSKnc1Z5mpGts83tou8gQxPFd7gKo68+vDa16O36eQKvyoW7kGiT
LOoh15FJ1FdCq1tPXVoSJYnjlkvnUqhvqtFjdjRVd5wOdPeIslIbE+nFwCpy7Dooea8U8iXlJmSl
rdzW7HNJd3f62mKZm4s82dBhVpIgfckLAq8Jcf2GcNqTBgmXjI9v1A2U5+YrtbC5Ko41ztKb8uXe
rMg5AvfoXU0ap2sShaPTxD9u8P7byIxPdyxTO6IC/qDOzdutBVrxH6FdoO1VnnqthLsWl6pXmLO9
EMsKiA9G0CWnwNyNWGYrRZKcPjEA1KkDkwbaC2krZtd8Dx7bGrySfbDc19vJhUGhZWnQcv7sF8Z4
Vec1ZTaRcnZtIYDlrQ4rXV6+W1S0A2IjU+703p2mmTNtWwjg0LrKXSYo50QLes36lV1avdDClDN9
5VvXxtTqrxmy8UEojHchh+gURShGsb6siITBMImXjf3lRW3KoU2t1XmgeFw6qFYWkXtCYfTl646i
O/6860g6AoeGIFGEw/j5d/kD1A+ZEQRjuHUofxtRBglWrhHyUB2RPofYrRHavGhWHKcpjILKYseW
Jv+QwkHKISkp5WMKAJ/UCEAduNWNKa/eeQyJ+mQKvEIXD2PRoyO19MwTLdG+7Rbp9IKGiuzDaIxB
Yy6rZj8zc91vml9AEBRk2lGBzI+YyXaUxvRTIofbmWQOpmYPtAre4Kw1STFupHT/443njVq88nOm
wzUhV7puJyMCGP3PsA7mnTpJU8N8o4cOwd3WcFhBFi4aXiIWfYrZaS+HDJ8cyn2Gj1x6MA51tWPY
JQ0A8XJrgXQB8HEczH2vYWuTch7/PMqN2Y0D/mVM/ayGfpEMQv92mxcuBqBDm8+xzHRkbrrJRtjP
i6ryswF2CqjyggPYTO+CNLhv/6IE869RZVK+yMMOphaG089SzW69kFo+Xuaql/VBM7xXP+92zeAW
xFOTZxHu0liHRVbOzTK04pOTf7v2PSFstrEIlM+yfr3r3GezcR/Reg76j72Sg3vDBlhzNEtTlBkS
0H4apBT23gxEexa5BM7pR6LAkjZdxi3sRFyjfiGtQs+9qt0EJE6Cyswt4MWMNF9gegHtp4KNEiQW
WWMnUEtb/SJ+sMdcK1g9nwCEw/yxM3OtKYPMCFEk9evemjepnWFbhBCW8eNH2slY+D4hAf881hKW
FDbJbQ1/ccUfrkQ4FSMZkVl9sWQWojmP/9QDFPlp+4Mee7aq7qfSkNhG/8esRfhINs0KIWusHwU4
2FhVP/8QtfdBjURbHbDonRFAarg3hm/AzdWJrK0TRqfuHpV0bU2ApZ8O2U0gYTxkU4WinkoWtxl+
kInit/dD1sAoNxq5FLglfjQsfpXsKrJ6LWh99ZbHzVEkYrexd5Ao3wX2JiayBFFJq0Mhy5IX96nV
tdlmcVixh73Yftlf0AVFUtSWLSGfAAwjZFRNlpqBamAGtm9RkiIXfzOnF5JeWG+4NDvNmY5KsHvl
onEgGah1ACl2DgvoCoepd5nu2dDENHa/3Qis3JNRTdwvuw28+sZsgGre2awxj3gsAppoOKhPILdq
bqirWIc+291jsRc7btWe39bCftZhXVjcsm8r36Mj/gqe5sj3rwzxTN7BOBl/H5K+5hJChLLsv4o6
BUE0e9CEkMi0OojDrlDZFqCLi1k92Y1Im+ZlMuj3CHaw9U1jmyWNxi2hlpLujlaUJuHsJb2xVAq0
O+L8+iE72o2l9pNpDUV6zzTTJ9Y+oju1eJhB1ia1s4ilvNI0huuHNRvju3lE+t6X1Ai5B4fSOU1i
Fz/EyU0ARw31yrT5thS0AZNMkMXdEL5hgrN9R+yrF5raXTdRCH9qyadgd26AQD/pPbOkyvZ12mC3
V9DwElXf10rAWw7/tDKaEyDWYD+AaUp+g59eJga0pLtNjPfEEjgVfB4pUZSrO3qw79Ly6m6DZDeq
oF1UT8mWRV+PSSJ2+dqwQhDQdkORwn7uDqvXir+/AzCiIajfqDn0/+FmWsI5P5jj0GdS5pnUm3ff
omKmgGI4oBYYPsNgWLOdnpe2/BHupS0aV9JwsHEpk+dHIQjfDFGaRc4ZGBeCaIlJCCYkyPpEiYSS
GjnhQRILynYX0wzeWjRNUGmcMA5/zFIYgCSvlDZaU5ADDc2PG57+/pvomq1gtUcas5vG7UHbj8xO
yASx51556iEeFllW2Zv2KDXwNxtDetk0aF9VEPQkhu/xqPFRniT7Efn0cYglc9dt1pzZ//6pBMl/
MHh1eqEdfc6kQkf79QlbOO1Sbu5FUq0lgzNVirfXLjUaKIqCNGaDnrNicJPOSCbEsEx1wYGnyO0D
5Zjxt/msUG05HdZaiVFj6L6RyYrggXeLd2e2jfek1QC6rNcVi12PYon3JIdugCD4nYDcUg9OSeA6
qfIKzKKTNRMPIr/sK6tGZmd2tbZonIMgJGsaFRYb3+NAYYIOZ54RNLeLlyJS1EF+83LwY/bpKwS0
62AFhtEydZ94G3yMa13fpp3LiXmK//pR57yeCQRjibZB59tP5gOgd1Bx747P/8mzYBp6HkDfu1Oc
mwEY8bDntheDwAq/Gi4/qfA3CAbzU1AjjX5C6cU3uYOhV4K9ueBvxcia8+fRDBZURvfopl9bQtj4
9AXtqN7JdKoCurWGm/cQJ98xdzz0ZVEZI3LxHFy/am6no2U4Z0YNfZPxulXPEYx0Btqg63NvPNLc
nNOJ+HpsEqIFkOuGLVl0bU2t2AnEbJVX+ZGEdU1EsAT2PuVNOCT+4GZUny06OqlmGqlzrAmvPJmV
1alYmaeMOi1tU/U1ww3FzjAPtFvqpNjnOKodj9ncrWuV/Hjh6O30Y4QAUIvMSHdUjuNEDgcWbtwr
crwzOElX40a5QjGOrI4m0ImLnMhkpoWLFabaRssqwlx7ZPxUvwpbQh5fBkTDEQx9dzm45+cYIUbj
VRIDe7+URjpLlSh+xkg3tTsLFYbHZy4Spm74AFKbxEcz+HaZ4L4BRpRKgnD3Rg4PsC4XKDTCZwPt
/Lnq1PBT3ncSGXhYSKq4Y/UKNEd1WtAdIzXGXAtxKwjuhzTNJgYUzz9yHJ46v2XAVh+FMiQaULKM
0KmLFOLirWzf+VNjIqj73OEMUpXJNepcObbOz8KmDAV4IrTJazjjEWzpTxOINovpe1S75JQTGkZp
77OerukA4MbzLP1eqcXSZ24taLp/WBKZ3QSSHanoHKA29Njpjv76tGDVXgks2tnE67Gm+JHmHACM
+5uqll/fJingjc1CS5RF77Zg/GZJ8QIotSF4xLaFoyq1vLSm6mYlTI85GQz32l/SLsRKTa8bbebh
LPJqSavHnIHxwipg9wYV8csYXIS7hvFXrb7UCrnpg98byObPpl4OCaBv6kRpTb+QX9JQ+OhPRsNG
U8LLHK1bREIuYnDVPfPvP2ahyNqJl7rTrD744XhfW+56+sPc6LPkmtuCIQCHuiBaoZPDT0mciaeK
HPOFMqr3BPwI4hHUNbxokzPYNGvZ9GKKKkTM+H05u7d7zlVyr/wq+4pEqN6iBN5ovcewPXnPY1gM
33tTAXrmdtFM+gKSK0uxS6qIHDFJH3ssoGxb7Bfo2X54ogGzHyM5wPMKOm+kP7vbZ5plxMyH6O+p
/O8c1jkB9IRTQ/drENUJXPZeE/7TkdPWYvjhXcYvj4STiA3TDbEIcuGYLWO33/xrnimYo1lBUkvP
23MuNMpyrlrOAxOaIEiD/M99n7wW9mZwhvjOlpfr9OVCetw35puTKfwX8r2GcN+Zex1S5ZlElh1E
r+I55zAFR7ryJQUu/pVdNJYGFYdrSqV6ugG8FqJhD8r6SUVMLhLBEaQHXtro+0q9D5yLEv2/pMvU
eu+6i3mv5WY0WsKkd9UCRF1vDAcOHCJiDw2znNmbvIZrbGp8GGzPeQSVrQgwCU5d9dbGeC1NhSWJ
kAn2Yw0m2mpOxdAOWoaTIT6NZWQv+3XRlARfjIlglYkzuI80gXtK/NpcUfiztzwXcAX4SgTlhC8X
YZX6UxuQA8IwjwEn8ji7ANWGw8WZy4P1F6qBVEDBZ0uLkbdo28fzKpqQeUSQhod7FOR7+UIkdwqc
8rUAC0plD5mdLuVnro5a60ERiswNlZNn6JseeulbjJDiRhcan5MDyrTszxokTC+eae3tWkTLRTg7
uUw3IHsGLNk519UVEJnJMn8h5lniLo1Ia4uTvVqpvqd0fTUK6hH8ATglNCWjZnPoWX9W0ppmVbTf
LrJBmnMiKdpRFA1epYlzVr8etOsxuFgDV4/FQMQT3TaZBsk2os/c9GEgSIaBAIchg4y/MXKuSEwH
89w9hCQ62SjBf2fQMbEMxdYi7LkcKra4AN+GBnDfcxT5UpmAB/cUMOpehw30jQ9FNu2ucRD5Cvbw
3SGcWlxSp2CMv2C3p0DYo2G561TwILFJN8Kzb3a6jEgcCVamNuiF/5TAm+GKzxmNfDjenslemHpB
8wdd+j1SIU04o+ngrv+lxIOSQWWkPZ8psq6PL1JHe14aR+9834s+QBGMHtNpDspfogJeFkWQ3XFI
MQQImrBdw8XtKgqgbLkAPNny0qJJNQ2y3tUzkqi2c7eiw3KxItZvqHhk8T8G1BOQZKSwzwVlcV5A
Hmjb0WPuA1FiLcQc1JW3AOSUxP5O6s9ieGCWZ3pHyrIJdQAHVSCkjSQUVvpCky2ZoZMnxZDJTgdL
EVuKKEHNkDuAgYzpnnGCbTbk33XZRsMmCiQ8uVmcET7KpDDujNQl8K6PjAeKpsc1llel96/bM4se
h9VAAY8L2kRR1VghuycE1rUOO3UX3HDlmvp+KfC2eoqGPPaz3Qw4+6rOtPh/vfrddp/6VC26qhbp
r0ERZxaXid5WVdyjgJtBk7IEzqRVRF7czwVfSE569ErNzf1k7Jt+vs+5rrWPEnX+AajNdUq3QDgi
E3QNhVZ/ipcaZ1PsvCT12ARoDZbDdjtFP8H8tdcSqPNKHtZiD1Io8BqRt8plIWPhy8Dzq1CZ08W/
DzD6HNsIoEWoQLswBsgiVKRhS7I1P8+sruOnF84oMP2G1jYBQmd+XrdqEjaeVSkxpnnL8ZYx2E82
zn9/dy8q1sD9YxPyK10RdAHa5j6KM3Jg1K6twukapNbc1J9SW6bIslbWCM2WALYpsuToRJWDhHdW
Fy6tYdL5sSNrHiuh5HawqR12+L67WGsmqGojosk4WU23Z9Ai1B/LyhrVNd/7971iDWxK+JFXtHMA
bGx1U2VG0k173NBLk8tueMoXqAh+27AIzl/d1RQGqi1JSnP9YGnNqEnQZptzVcfaMKjfEqu8MXGT
YRqOhtH6eMW5tHwEvM2rd8++iW72XX2/kwMLc3j+gv5/UL9NoeX4d/GQVFE8ktsJAi1fUo9QldgS
ThuNhNP4Cuj4IH6DM0RpssvAbL3Tyh+UOrVwo/aEpYLbl7Sj0SKGVJ+runQnu/0iA40Oio6T2j9f
Bps08SmNtnxlKwU3UMX/BXQyUu8ehlDwX2Jr62ng+07lsQn8MdLa5tVPl0uqN7FUroZJy5wNeSy/
caSoaA1wiPHvrPZZg6zxQNoBPC7A0H5xIlFDqy4qcM3EvwZC7uIC0W123E9h3jFS1KkyZdAMKOpn
gK9D0IcYddYKOPXr7Z8SLTUT2MNrDDE6jEqChHq8rhO84KHdZeeVm0FZN1LQINwKsg5BIIkWdsag
vylcG99KetQtHbazGAr4b6G7WzOdXhbep7oJrCZlfnF6nx9k4lfPCajSlFOd2I4wk6ZojIkgoSw0
M4NuNYOCoGdqSl+IreV57evfZdV/jVnJcEq+iPd0E+oQcshVkEOpknWm5+z7pj0i5EvZzhd8v1rm
J4pph1/mQTrWGxiZrz1dNvnICAlS9PUJkkYgF+YrPGbOgWGQs2tu1aSeWoNtLuMZzbZ0nJ/1D1Rd
RhNb1ZWtJbPX5gUzdh8RXybs7X/DafDZG0nQOuhaJOeMzoZ/e8n6OQQk3u6XBcPeTC1lOhHS5aCo
Weo+72ZEqdWPQXxIbWZm0VGBDuzsWW9pct7lRfyUwOSJKUsvF6Zz+fzfffyqRQ3Ayz6ZJeHnaa0J
CRHj9S92i2RMgRbao+xOV8Dq0AX0Hi0EgZmxGfRTvu2Vo6+jWNeOP5tv86vfT9WbW0nCl5Z9Ngz4
Ns95edVV1F6dUe3AsUs0yEufkAwfNInS5Dm3PkPJ6UzeyGkxpqtY0D96gAW0i0EE+09Xb8L21ij4
u3CWeAk6KERZibafkqQEzIgibEjO3qZx7zHLsl9vq7yDLJj10rHy5fQJ7Ul30tQx/uhhFfAuPlHj
xJvMH9708K8/hsb0czTsZTOlGq2mTTpA4pGQ6Wfi5cf4q2P9O5D66B/0zV2w7Yzc2hfBBXBnh5xm
sfo2GHuk1ND0x1GfTc1sNE2cH9tYkTJQvqrg4CIZpMPmer6v4LNAhSB13H+LV9uCSE0alXPyA0wk
1VY5HCevOHYVmg8IB0NQgvm+G/EfpnnGbXnMiNoxU8dL9DcjYFpkH67pIJpJtFDv6k2QUd2PuM0V
HYGZE4f3WWLVIfvjX4JUzSBsLKdREMOpEC4u30uhCc3CdkrizfjiJgrXh13qgKwXgCLL60oBWEMg
kFKg9XHeAQjNu9Yi5Ligh83q1G4EgM+bBcD9kcb3CWh0rZQUSABaxZYEWNl3eqmakndVdXviFNhG
K3cm5UUY8SzJ2W2EKwH81zQfQSfxBbguz15nCxXoRpG3QWDoWUUnf8+gUN9G7sS0KEfIZrZS21p3
gah1/MVYlG8EG/M7PxZCJgU3FJCyJIyB+MnMELXUYxqwQrE382ofDUQHYi+wJ8fmMSbIV6otJPg7
pcNfZs6DuwRWIm1Yg2m6djvAuVgsEOrmT7rhgYIqASchPUE9C/1/AQwLm4uD2vhfDcq1H4xxclsr
fVpGCvg9hP0068T3GpHBzRrnm044U7h0jv3QrKeA4kaExQvAqtjErsL3a0Q62xkRbltSw45TdfbM
3JoMEl9Hqfpgrwg91lzv5HAuoajtudRczZiBn/GUEcYj2m/GjZc3L6kbGZw3rLDn+TDWicW0Pfhj
fRwUk9grWQqO+/Uzqht9PU+4PtTGhrdiZWY+ImOrloBNnpvsGM91CQGQtIxeTRqmx6cfzUW9LrFu
SbEnqEwY2K41Oc3lo6vo8HJqGBVqO6S5KITQ6/7E6/JbQ+H8kxTkKaePQSt5ZEnTXSkI4fxz1nR2
NxA4gsBDXnV72XSRUsKQbmez1LDE5GlqceThBUxnhOxKIChcJjCwy3/FQWsc4gvWoI/hB75nkomS
/Fo3XaRmWLtUKShTdLF275DXzyi4GaNQip+nWJcpP7Beu9bFQJn55+jPjihiyqqav26yyYuleKNu
CSxFzECi2p3S8Y+sdwaxnVZqK+7T7pNEANYfvcA4M++Bgn8cofgjxla3ug+wI7x6WSpv6AotiXY7
jukBya8HIx6C4SoUQbbsB1h0lgw1jGXFZgxvK2nzdnk2NphsI58kqa7DyiGZzaB+GhHKCQS9Q4Xw
Wlif8Ywl4OhqDd0hMJGaj1n1yfVzhi7dmEIpoykGI2lKOF/LJabjat3ydnZuBOQNcy9x3zI6rshX
hPj+73R9bbeG2S9vTjnw03vexy9RHfdccwvGPgCp3XjiijeHs7BOmeWoZVERHUYD76UA1ZAk6Rr2
sAnU57WJ7Y1pSWcliPXw6BzFv9fpJ8sg1xMEJl8rk5ErC4DCDdg5uKIXIdlEe494WqtTfGry3QYp
tMgyO5PRBx3ZM8MmR3y91BjZ5IWKDMdzBbeF8z2b3c4BU2PkVoGgVu7VsoQahCFyRNuxt8Wvp4KT
JEjodZ0c05yHmwc4MIi5Y6O61EjD2mP/py72vzdeY3TKvXAeJQwVF4lglj9Jt/1TED3DW3TqH1gR
wlELW1SHziEzRKYopiWZKbgf9rir36gTYpq61FxLNOj/6bnS4Ks+w94RhIYzejkDRpmnU3Lkr/b5
8aWMExpfpRk6Z+bqXcOakCGowPimauUwp583mRlB0qkYlC2AnPr3ZW1j9xXJS9J4PmbVmHiDSabb
JWgsG8t1BSrtE48QbBw8U2Lo/zkaj3J10tX2s8yl6MWfUoqjEZKNyACp2seyHpfBnRmYzqq2W+Ge
DgW6QHn+m6T0cmKynSx37978Wnv4jPhjZgfuzVw5TCgtybKZYlm7JyHFC3Jixhtzm3U5SMnfZBS+
oiJl4bZ9HopEmcWF+kcZKLBVDnpbbBlcWE4pvaEN9OiB/4GXo57jwViR0vVsJU0KAp67/Z961mw3
m1V3CLiBeyZG7fWxdO6dUTeHDKoJK1ogdpMPcYb6UctA+ozia/sgwhUbw96MdNTzmJR3VcWQyA/H
uAtZpnvCbCOOfyB713wVMAdzj+FXI8yOWCc0X9viZEptW4xdDwRG4pEuJBS7kBQ1fzwSbeEBS84l
AID8k+5cJ0CGnNL/zE527eRtgpvIb6EP0b+524lLN6tWW2M+cbHDnM13Q1l2lN2SisRxzmxbGKzq
WR4/bacAqbOA1sdoPpamjneHLVM7/uyVp6TUjvXPs1hHEE+OvR6wfl769nTm/73AG7r0hKLhStxY
R0diHHDBfW3eOm28FNkJKu7PoghujDc5MsNTzsE3Gnj6vLDR1Iv8paEAOVoAj+N1T7uqCfgurytH
f4QPdluMqL+PBmwlezWSeg2rKGmeSrXqfsAGSRrGxniBa0vMuBwVaQQOC3cWPi08zPfDuzcZb2Rj
QUx2GiHT/pUd2BOZUvvfJKijz4jpwCzwWA3yQEaKeH+m7rXxTFbIuJ2eWRSJlyHf7ik3Xr+dAlir
S0uYq2vn0/zPusXYA9KFmJq+QjHnthWGD4UtTvOwC1fUDqxiuq1vnq7T7KODtV3nC4LfPR/6sC6Q
lDf9MIIXmU2cQKpIk4WSeD2Vb2TGLulIxtDVkFTrBxYMruSHBc3rkInTqzXrSK5rVG8ft34S/V1D
SXjnptmoyY5ydrLPWJ4hxXs/WEGaS7XdoS3YTT608TggjJuPyqGz94nDVO3CtH/79fmvM1Xf8OBP
YcbObLq24yGWxPBugURPd1CYEmOIQomz4hfJt/iKo6XaOgxGRifuzbl2m3wKiD/OXgWUDEogBVFZ
fEsQ5Li+SdNXUr6v+0sKCocV6JRLp/wa5jO3CgHa2aC8czFBLC/JGlPd+ToxOVjAUlAxr2HjplDA
iZmRwRXtu1hHl0u3BbrvzaKc9LYkvh0VyhOd0kpbCsfP5QxgpmSsjzZ4dzD3CI97LU7P4wfNkp37
3pJfbOkdYIJg3de9DTgdvy7EPHpKTDRzM2ANsD4wZGZ3i8M2th/ei4gdHersXe0c7cjHjG6Q7Up3
CBuTwuTlxBTftZXSLwMyNugue66xOMJGk+EHXGJprBegiPDIFGxOWxeqH3h/uTCbmZdqt4U64nd/
y8zd5AzDgSyH1PBGQIsBaWPnhVsh5e3TcO3TyCT9ZyD37ZZIL8xI4Ftev+x5PmEsqBVEVAh2fuzt
5lvYTh5o2gPbA0kK499EvGd2AE0300IVl8sbHiTZEiPKwa4yJH0cgMIbNuS+Ckr+LeK4Mia3MM9w
s0reJDdLu3J8OcHxQAvpdJbEmTuKV6a4+qd71XTEvg74epdoT2lZ2v51cQKrwXkuYHjb1kVW8eJH
QjOaZNApbEzYuBnXvqkR3Py2jb8lFCsyiiBN5RyL94kFP6Ems+Bk30QvJRhR+a7AYu5/Tpa1gwu5
6ndGXj0N+NzEr4Zvu3meqaqIsR0XR7+XxbQxUkAgkpZpHHIeqITqDveA/qQU7ejPC5hNg65EYkKs
XfqVPEP2gWC060XR0f4O9h3B4ia4z1Z9dV0yP9toGWQr9E8X/uh92IUvxufDafrwSjgZKI6aiyai
C29gwZNzL6qBEumZHc5HoMGYA7qtVUgK7HoAGK08A4XvYolDFP4YoY1De+haeA3kRmO1ljc2XOed
K+/ua89C8NOS52gNVOx6z2gRWH0miD07U//zveg4XHJ6nyqR38GfssD3DZvlCNHe97f4WmhGALw7
meDUFwboBZtfIKmw9bMMVYx/VHm5BL6Eo43QaS0tcAO4wNgQjKf9hUe6cyuZjOpjxc6luyCY2l9x
z7x2GBpLe4HoGULtd9B/ZxxYQKuBcoSfJRa/aXZXZ7Uo9iqoLNsu6QFFUADpdkd8AkQqcIYcQiwh
g56wLzs/fteIma2D40hqBU0cCBaCwiErZCdEU2x9RwQ7pgO93JQCDsrGF2wkoVReXKoHbo4SzvrO
jmnCSi/4JN8PRf8VoB72PAbZtD7xx6KGwxk3L1C0TZViyGQBvBbPR337DuekR6AlLdBqREeySEYr
5Agiax/lA18mAUGdQb4EjOxQFqMQTpFo8AQES9TTuDg7t8c2Q4WDd+tvhjV7Ikf3Yl+MHZW6Ha9U
yGpspSM9Cb0dl98K/2RK+0JGT6605PCMDprOu+q/903taTZDJ03B4hLeC0HL0e8/kcpWM+6SKUgk
HOoc5hZ47evunPmpJLghpH7XPqEhqpK+6+SXO8DB3foZBQNZJyL4WzRoxejpY4o/UC0fJn3cLJ4Z
Y6Sqgda+xwqtEmzocBbEQurfIaYBwe2V4wJ34AbGDWKk1v562hNd7d5AdPbTcJK9ZLc21vNnFzTs
qPRTFIpfAtVGQkR0Y+HfsjIVpckd2jLRzaDtiyT+HXXZ/RaXWZ0bRJkiMv/nJQs4ZTPcuRJmyFVN
1e7QYu0gZ+LVwSFUyBzjrBrVc861r70dD/QTIWOm+Hu/yxXMilxbGk5ltEH6Qlo/GwMTWEdLpaEw
p0pNrDNOz3aGbx6vHK1uR71mtAjyy9dQfF36HUgSU7/ntmJ3Jnb4obJhRoxNvSmhf/aidZInczWl
A6q731QZnj7QGgqOPg5vWJ+/ypIzQutHuvimCkia4uZsLYLgoBnL6pGqkHWmbq5zPOGBnOo68Pib
VPyn3FKC/q1CRZZPhAesXn85YJJmkibr4v9tnhLXhh4wYI85JM9fGUtXWeZGsQMbMZixMbo+F5m0
4qMsSrfH1T3MTngg3q+nKDotpePF1nU3d0/PgMV03Qwnh+NTTkEps4OQOVq/N97CctvdRKw8GuIb
5izgP0j+V5vpKFDk4kkaXvoTY70UchsKiLGaL9VRYLuCvsZpH2ywAElPvedIM/6tAO5+SgUw+obI
A7ks3aVqSCQgQEWkmQtyUr9hiZtwgVh+uFeYleOfWvspwQh+F/Nay7huYpjWN63lwQinjlOyDeIb
wcZk+QHbZ9as3EvALHHl1jt2++gYTrZ/3zKPAMrvWJS9+adBcitXFPG2ZsWytI6xMWm9OTzcbZ5j
AwtG+5n4DkiHKo3CMxNQxU4CZrXscccoCsoMDzh2knjGQJPKC2hCDqNO5B5ZnLFKMx0TxGB55r6Q
vbVugD+6k45Yh3Lg+IhvWgCy+ryO0RspVO2D0bKxMEOFFlDxIhU54anUENAExaKhBi9GRd87lzMp
TE0kHQTYIGiwNRrx6g8ypWiDtfO9JeyuuabWfZOUs7Mlyiml2EFCzgDqwblAezDp3kuTyCK2h6Y2
lH3yN/foLi+Y7hFVER0Ee7ybDUM23EY/Pa4/19qG+qnUnuXodySh1xgi3GunCCEG7PMx9MfCgtnM
lT6AxY09VhjkZUs+wXkPrUI5e3v1LPZLAvGMXMQipceGk1DZis7BftufJM06raYnC0UVHKKiGjSv
lWWRhEJzfqms/lRaDBM5S3wLpHF1BSUMXmO5Hy/FT99WdRlhl1TZIISSpbOC8SSvcquuGbHH49eb
c/mdN4iuEObbcgqQUJEd83N+hF1xc4Bk+ORugHCHpWO8JhF8tdkOe+bXhvzXqxfUZC8fwD/P0pmL
6WqXvTQ9/WKK2YWd4Y2pNz6uBJnR3btW87BOIj73BvM5MZCS1FAeu9Gyv5V5gNWQMxHCDdOLQA7e
cBmdgV+18rZpPNzYtxe/UlHm4gPhrH4fO9VLEjdMG4bkoTWjcjC7vQ0rMcx2eGM0jM63q1MUbjSl
EpY5RimrreorOVcQxq05eWxNMRT5aO5O9Pj8aUjOjc9Rp0uK7MCQnBgzdYPYnhNSdPl4f4zVgo+R
ncUaVsGvydI9xiRNlk/HqLGQlKyGpKNT8NguPLU8aXd7xhL+LM0Vt6WVbW2VpBJLbN474KploWW+
0NONeFnEqx1pFltSmz2wjMIMM4oGmTj9HqJqd8Cggq6zl4eqlDUphBUonrPmbei/UYWBNj/1Bjph
I6VosQNwT+7VN0/cpsnbJ7HcRLwvpuMsaLvTgPCJUDDFnimYi1tg9h3V1Gs8LJId1Yg2bL6LdKbw
lIO2MNMHH8m/70gAO0vqtBnXnVFpyHFG8csEb6h6Uygptt1elEdtOZYlOVozX9fipcxJ3uCJtMzB
jZw9CwL2syLTDnnMGlDvAdpEle3Khh7vrlw2GYFGLIqbKZtOi2ZeZghPq3eWvCB2KdfnYeFpF1gh
fKw1D/PYbq2HKXWkMif+Kjcc9nqpglJSuJZ055ozsX90Gz2woImEX4nhXb2+qT/A3BEOYPS+suDI
xYyKV57m/1uIEWHQFwyoIBGzGc3HdFiO2BdejeY3XzesylTC2X4Zh184gTHLIl5mOhZoOALhHhzx
JUfGzR9f6ICTJGuDNBBRDdExlElWzHTf9NjeHO+EODpm8CWmAnRhdqCPxynw1UxP3+sna2BoD0Io
lWY5wI2lZmtf9TCNruiSRa5Osk1tp3r4Wl4GEJ0HvhZVNnuwK7R8ynPGyL9TyAIoZGrg2VIBfcbu
09na94AgmaRMO2odb3tV50GDFScL+YY8QGyq/m8ijDe+KSiOvWZOVSw/TmwTxePE0XuxftmnBgR1
2OC/H8evWZbbhkpdI7dmMXDj0UaPSz5M2vbpwYUrS1rwqeZhs5vXhV87sOvo+jh0bEvu25Q7/hMz
KeEorCp21STa+9OQRbIHouDM+Ml62yRZXO/z5LjkQeljY8tqQYsGj42l0NszOayx8jAkhpVySAt1
ddEgBVRVa0Zt70Tr4ZK/MqeHwnilJevqb4nffX+dfXK6vNbz+VExD+NTwDT7R2fVzIiGJo4SmXlW
nlUKhVcMxbATRX58T3uSy1rNDXeLAR1ulPbyHmQ9IqO/RPx+5/6JamWTCRNL56jXWnwez/wI6l1Q
JOdUp7TYv1+bCUHIF3B1XizXoC4DDRjigEERtPeduQnp6emgDqUfqj7c/ZK9W64bW4ypXpEbPG9y
Sdt5/FtW4z+OLVZvkPewJpROEc+di86XTCrnQlAPwbHwebnaKkMj7tZ46OqHP8QZohJEpk5tYrUI
Ir+OaxGXfLewcu0AWn6zP5vrOq7VkWWoExh6kvRNLJRxw9SWypY1hshMsCZbLIYjTbTJPLhdn6dP
8J33omWlBC4SoQo5uen7YjhcqTS5oI1tOgv11mTAiuXqhifnoerB+wLdmMBKUQdbP6RzPiFSvE67
q5iZq5Yo6Mhh8n1F0kSYDVlkCc3GexAd922lVYdXgR5m7cgFX0jJE/hszZp4R5wWvEtVgap2kSE3
ZOpLQCkkkXEWMYrOYOwDgCGf1mP7UHeyT6gFaM6HYfDie5mD9cvofJ4dBOUThPFzhA5UVYEHvpAJ
i2VmqbEiQN/pdJ5CO/+ByiQ5fkmupo12iy7ihmhkqVZhrKYkFF6uNhqo+ypAIaTgCceCAKsbwKAm
/TZyuFj33+rCvGhRLFrUtbKktRKRnKAC+yinN7/ewEz4QWh4iHiX/qUAufOEMB6mkgK46VGQ87nH
jHcdP/PU1umsivg0X//udvY2TFHWP7r3PURCxBYBe5L1Ah4aOHmQlhVvHBk7wmgEzpk1BbJegEGW
AhG28x44P3yZ9duUZ50q4w5pZyzHVvxhRRbNHFNg+H37fGz8ILBGVPPruD47wvkupwmiLQn+YFUQ
Bjaqx6nmriIq5K8z+QtShccd1XskwAzstmEjqwZPwSrjVFYG23KfMzY0a5OlsbF3armr1arYDG5S
Zoyva3Mc3/tkhJ5lWsU4a881PMvBkMBJ4FEa5R8wMzUuNEonBUhpss2Kyv0u42shI0dFGH99J4hq
9x78DrJGBiqkczq+0qBXUuJuEwHDx/8a7qwRThbXfJnvMweSPZqgZeU88wPDScH89C7eoHdmrhx+
kLJhLAjj7c1Kiguf2wRAULzEZ563XP8nl1ZcN7KzlgeE46/a6vdD1Mqwf1xarhwQ2jyEstmFwckK
34yFAhDVRKk8KusxeeDH1r0dJQd+1TlSj59N2RJWE/qROlwlegJqudqQhK/oW94GzgA4vBHDp1aj
ub8DYocDAXINMA8nd3qLd1bUTRQ+LItRmOJHQqF8wAScnhkk3dtjTS8wq1Ce7Oeua19jluF31jyp
5P7e/e3S0lw+ZQXGWDKF6udJBTHZjTxSwbf1AbSKLpMfN4kIjAwb1G02B3WFGt+CA6xspBmapb3d
6ub3AH2vcJjvSRerp0XV0ioIXEjqztyiSKp8tg8TaeWgnkQQfYpsSEH73dxDZVNdVh1CJVvxFXez
oUyxYfv0oPHimvmGAcsbX90GnmfXr+FVIo+lTf3hHf021J7W6GosA0g51s0Cgq7jYWf6RWJr6/e3
D1p/IaOm4fA2PRUpCw89TfnydYoQ4PIJOt6jvGMwYL2rRvG62UuvfN0JlrYY3ONNxsW/xFqy5wSc
rQ824rO0twQHG+g0utKJ3REdniZbZdzHS3eXMHelOKIeEVYAxlJFQHra6GRBBr99kK+/V4j5OG94
Zm3UAhD6eqeTLHW7SF971qkRxjOmXwvGv89sFn0+zIzBL22hIq1arEGVNhqyAvWWFXyDtU1i/onW
T9qaCBswzopnQ7c3xcZ/Lop3ZyA6kJpDa2MP8Yhgyi5R9E42MLEx4krlNxSqVersGb+PsagNbjEe
ddDekaAEjXaGkjrDO9dySQQDYW5KebAT5iX0CrhqQsH1c2SiP4h7O5lJ4DdSmduBnhMR6gKqHlKx
mrEg3BgvVUvBJdW5XIHu1JQZixU3181C69P9rGAv3x65DLwrTEEZlW199IJrwNQB2kxy5Ip6sdlZ
QD/wKU6aARXEQMjPpgDySIQhqhE5RxbkZjeNfY5Ws2tOcb6QXca4no34vwj9hT1AxHn4n3rl72f0
A3ZFEenv2pRUq4aRy1SanCMFsqpdPhWLlFfQq4c8pDDvkNyJL2tNDK6ugXjjVD1zF91b4ziv5zdT
Ek1ZJ1fj0NgNv7U5YBCGetIgWVl+FTxYnYIMHiSX492qOT9jkLx5VTgrrCM2rGt6x4/U/OgPKaZZ
I3ZNBOT1nKSUbMZ1itm05oOWDKF95L6h7uUnyvaixzZJZkZDzjwF3qUgObLFE4pHzSzLnjzZcM0t
PL2JWCVFDc/rCEo/2VrOn5VP3BjJsV+VQcvyRJ/2j2qyZW69qJm8EPkHekdCNhM6/1utv5JplHsr
SQkr15iWHC79TYQ2Aqazo00vNg2Wujnkia7C/SETPxDze+DlRemCficD8GWCoZCUz/SBV/8zP4aL
ZYifScsIYeM7YOAONztA7F+0ujKCCYufbEyaxOU3OM9W+9A/X/C3F3OoroIYZ4mivcdiXz+1KRze
3MfkuE/WPUtzylvNtKB1PDn5ULpCRYvQYEoW41x1KYwZOT8ug6/ZuRjYQibVTOTkLDCsMO5RfDmV
fEMNr06VZbzAT28nbB8NOU+6lA7sTmcjufy8in9lkMmZ46qQKFyZAv4Nd4T5cELtV0J6k7PD238/
P7F9lEaWQTx8kKyuisR9GDJ0+IwcsObf8hpUz2rPeT4G+0VYqfa+4swg6hCG0qqko8xp2uMrUdLe
z6xNeDdJCU27xBVqmx9Y1J42xzZTQX6kwcnINljsPV5XiHo+u55dAHZAz7EyCeOyDtSUd1Jo4tbI
euVv+pOCmxrk6JljpXjXG8cDtcpxItgujEdOHMNYAnFnkqq8g+3yLH1qEARS0RwNJXAfAWtwiObQ
habzaAdJTMuVzNyrHhNxOEG00XkKTcYTKOmD0O9QaHEjiJ7hGWLJVMp79G46cp2zy1YXmwgsghoZ
SczUkxo0ERqkOcW4rU5ldEzDDsuW2USO3OdRHh4GeomfWz0Mf1Jw+ERqFrRCtDfWwheChDt0gvzt
XNraQDq7oco/hbCQ2aIoj3F0LB1hBHoCb13ZUWZXAsL7Zne4maG/N6VP1mDoHaYwODtamCwhMmlV
gZgjLXoibjrKlQyBBvNhPES1G3CkpWWtvr9SJ0Fy3kid0vLZeOSnPc1x6in4a8l2nip6AYyax/ij
EzXYO/pmIm5VifiKzQ8g/CJGpbe+qHAXA3vU9QOkFZPY89Zpa/TAG7r3WTf1MieyYhihOgnkMD2e
2EdOdUoG86/jnuwGjGzbKRM9cMhKhb76nmZ5sORgIJdt3SphtCO1KVzOH+KXkaLihpo+ePh4MeRg
107KU43q2qclKvXIQTBmIVHIJ4TiO9g2NYykUZZzLstseoZAxa1FeH2A5dp+bqdIRV+hObUqHg5T
VlR7nZYAKoDVa0KpBb9gbYWicxuYAQa1DBcbiuMB5W/7R1rr5EcyXTDXQ47j1MOdb4UgNnGu/FQH
uOSWLHPdr2vgWFKIVwq8DZ0SO9G/tMhLnWuoq2CiaO1WlaLcEv4xGNck4Kc/1EKL01jH2y8wuIod
H74LfFQjGGsi76EAXMkiXb4P6UGXD2S95gRU4QTo7aPg27mgSkEOfbW438GFB+Ri08V6CqsW7mQx
ZJaxIVYKcY3HHrAxhRAuua5kE7D7KWgvGJ7PzAObmHhrWq5ci9hV0ifO4aRgXN9O9Vaua+MIXw3R
NbbDQISoJuA6hA424Zn+kG2KkzJ+oiWL3TCRlhII0Ay3tFLsO0RPxsXZFozg5HZQuese1kxLzLcO
DJIWbM4mIdBCm9NnhXxvhhibeJZpJfx7tZVEs+4imMdhv+IR9FoRAW1M5oEMaidtshq7xrfCz8V0
O/mRES2585Yolm16in6ReuHMJm3tOWMyn59/VjlZNbpLwyDAt1oE6tr656WBvUGckZQH8mpPPWVZ
ULGFH9F77jk81BHF/CMMWp4EFia+JiG7DrwHMnymEPDl2BFB+Uih9bL/vFQG/Jg08o/LWklQ4LIR
UqlTWSClTVfccrsHdbwD9NE0EnIMH5N/Qyz0yzFw11IPIoU2CTqM2pPN4eAiiKPtuzaQT/gH541u
TngPGhtBnNEMQZ/BhlUQgQ870urKPECgEgxTKZQbA6Ji+QuJkt5Wyr+LwU9slpTHOOhJ7q8E1hKr
PS5AMZ7LPgHVA8CCIEpSQkpdfpP9kB/LeT0VmMg73SHRGEXRcsfZ4o6pVoykRDiRScfHi+yhr6qR
3/JsO9jMUiraerpaj7x0w57HK+mWBC2op+jFoJ0mJWHi/0zHwGZ8dnvrgJATuknUan1lUv/BsOjI
OaU+F9keQtytvWuhjwTn1tZ/N06UE5/liPKB0mXi0vu7Wf3AJ/B0Kv8vKJPjI8n9QRFjftjtnJCP
t7Ohd8RbFGNTb0c6SG4fIoqIKYeNWGCGuYWnUBSrEwl++aSgITOOk++OPkQ3cnAFK4UVgsxVHDGN
On47rlojzqAYvY9rXX4vYCMTkiJ1cqx1VahQ0zPhXo5UgVqSOGt/t3++s1HRc8W9V+7mvcK9QEP5
KDZq9WZ0NRjs7TUXQDReQk01Fu9A5kkux8zk+AzlCvrhN+r7bhPOFIYoJiJ4mij3J3Yx1YJH+N+z
M7X55zqD4O+6HQwTZ39Xmjr49IgTY9739J2SfIp9MjY0uFHF0/x8S+eGmSAoAKi1A5GdPcvbUBeD
5+A5nhroN9eZyTYFgpCKDFSpv39h180KWmu3vwk5EWOUnAFxT74AYagt4bPgr9ASDRPrlo2rSdGr
mkT266/IgIypZ0YrhvMgqwibsKra+GL5m8mJ/Q3WiYpHTcsFnfXij8w8BOjCnysN3Z7aGW8G3orc
pU5b53ZIfJJun4j3DZ0E67cGZ2CZbwq0RPuHCJSCitEQFYxilcC9jNuQgE3n1ielFEb+d5pnihSX
sqjPfoRs1EQiT1euBA1WKgWHcYMnt5CQNlF0gIBEr4yM9FHI63MjoqlI0qJyzYZyPDzY2wJzk2iM
sq5PwEI1QTw5bq5tkV9M5c4Zi1KXm10pgTkGKwITiNCGFsZcwBLpCwa9nIyNcP2ysmYCwJrO5O8G
cOeZ83XhybsUYBS62s6FQ8IMQRwMljVYSjz7gd7qKn2gl9gzlPq2Oardxg/o7A8U5nWUFiY8yhFw
wnYkMoWd63eDhJHEJEM13Dj5XZ/KNjwP+ebLnNtUNmWQa6JAat8Jy6awrHEDeh3o8NBr6VAODrU4
gVoaXPFS461UXfSroAVy8YHB+GpRAy2Wnp1YDVzMRCY7gsm5pzIybjrYPkptrG+uXctTushWCh+y
pFoMPZew/5gOLimWYIFC3/GkjYIBvyanBt2pWzKf3bY4lswLiiLYGMawbsvEQqajPO606IPrIdtA
OzpWyK9SpAk0/D0N6v+6bREZCg/HiUNu1hDSW8w2NBpz51Ty66lvpLzNWf40+GznLzEx+DJOqs+M
Qb8KZw8NBihVkIfPk9vTRYvTf/oW1qEQ4Aq8oW6m50KqF14rYf+n2qmr0MdFtc1xwhL+xR1o8EDY
79ahSMQvvvrsk641rfyp73HiQZ7Ly+ajov+TtUZiq9Qz1F629Id+BzjFo6ZmjQ3V+XuxUgR9ZkQk
ELxfwvKa9icWkogKgGGuaEfmYDZ3dYO5ouUEmY/nf8YXpKBNTG3usbAOCN6XWSUOKawOVQPhMvnT
UldZnbRtXIOVPX2+KDsDeevJM0cKXAg+jX9lxM97BLMjUo7RyUKFYpL3IQhs5zn81mCFfARe415a
A4W8lwsJGhh6haOTKH/MSGQ/3HXZlpLsehXbyVXS+cgVuKZ4sLvXUX616Fv5Tw5Ck2ALmR6yikON
5ehWNrjIcYfvAcpM65D7eWhGWgX8Gini+9nunyVI1xxNQbFEvtl6iBJTh/AtX4IpuBGnWrO3J//V
Jpv3rjXnKT/qeopa+rAPUG3iNGBN0Y9h/K4sju3DMeI/nJK7JY22JplN3YtZgFmMrWW3E2PUnztd
FmjNZULWO48bR6qxW8qOhwWF2YynVClWdCqGqbBdgjdNcad0VqRAlWwAzgVBJP4J9CVcGbp4rv8q
P9hvk7ItpuZZmWd4E+29jV+vh/+yOAZeKTkId8w71+p70E8TC0MSQT1Iypx4ZhJIeL9HlBMX1KhI
/OhJHHnDWelIryJzAwkbpmmcyUAVMynKGTYrHmQlnGaozesJjAtRrtfgc4j8Jc0PH+EYfGVN0ygW
kcVlPMpHWm9hMXI7bUjgRKkveWeP6Y3oa5ikgvYVbsPPmp1hnJTlgDF93+Z9iH8+2j6ZButPzyOR
8OaMMDI7aDReEc/nYk0KhPt0oYMZAox6J8L6ZsYMvjE1nrhVIX8nePSUN+ohVoChVaw8JurlBBok
17urPnXhLrf+UQsAgxZfDpEM5o25Dz8kBxMZaquyFAByPZlCL4Pja2uw2A/fVeH7tO+4UoP5hr+r
LZGIxxtaqLRaGqjHwsVzTZttjgwCQW/8LCWF7dyNpetze3nn9GiETbx3l54XeebOfJOSbgrvJPKd
1EYB/xiFNQ6rqOa23uuUuenyeY+qzDZ+eV1f6i9MB1xjx/N7M2IMhc06swFynM2BsWcTpzKU0BgP
D/rn/VTmfypVhJL2rNE9axRnQusFTk7/Ld3uB4T/gLo8IWqQcdr2TXWdH/QpsYCXB8ZTCmKiP3dO
NsTBvvNEzLn9hAjjhxRHfBy0MAaAI/R1dPycCyXKa33lCAcg5TVM+q/Wo6skNdGrIJEaSZrltlrG
V6zqdgki9zr0MXXrbsP+Fd2wvAQsaadZwh0VZVSXM/dgsYiXemMpQPEZtCpxCHeUI9f3hTq1LrPg
JwgTmJNY9cWupuFC57YBZoDOsGZmlUJjSp2R8deoWe6uM6KYJ9s9eIrG65bt6ybTLZHcYEAmiijh
1jQJKGy6usfBuveSkQdlBehQa+GW8FVCg4ryLMaNxwfn4L9VZLH1dgdGtMzgF1Wn6B/VlpTM3wWe
uPrmgnha2yaUs5Qyy5WwIB58bTeK5yIJAq3EhOXPgnM8g5zXW7tNVQRR8umnz+zFNXiv8ruSOsQv
E65HWyPs3OoGQyyHsNKEtxmmp6qTMnCKUGK5A645qe0aaCqPj2IrWZ3A5ouYeAXWvTPqf//iA52k
y14ZDLAhN0Hhk05C2mo88rTiiQh9mVdqvngxBmpvAqjbOMMHZUR/L/MWJva6hwNGn6Dvc4bN5zcJ
ThJLCH94QxJ/kJo+iEyivz4TJXXe1UrI1YaBgb/O+feR63KSWwT4CpjIr9Z9Dtl50D8KsJr6ciZT
PnV6M6uvn8n8qfSdsI6sgXPZgS057ayMNDOjBRNOa6Zb/CG2JnEMudR1WhLbo5rWCXmZMwg4qfa8
fzEerdHqTYQoYonVmzz3lQ1FCA/uK+AoxGOet3TU8V1Jg26mjbzm4TH/AWrJ7OtrOHPJK20Fr0B1
7DS1E0i5mJK2c+lBSzDlM7wLuyREQAROfpO0IIOwuxesCo9NW9qXysokDdA9cFHixcEyCOIswwr9
cz2hYNfkbkG+hjc2Dysr7EHT/NQj4etAzYguO1u4GVgILG9mJS5d7PBmcjUFAl/f2mgAX1v+CMZP
1uxEFtZOqG3W7B9YPD2N5nPjpqySPy191WI/kSSssZA9ZtAtbFikaLJKrAibra5qhlckprdPB14h
TP0cltGiGYw9PbJRP3mWnPaUcDyKvZLh2HLUtZW4CSGNLVTCRvgHbSWCtyVTWWqTDyIPInue2n4k
lY+gZkFsiZqnWmwjYcFMJKCyUS0+3s+o0r4MevBYigeoai4eVIBw9hSqLFAH0eoIpxufT6T+mwMs
CtLnJTHeffVP75i2rlvogHcLuhTazAMASSzPNiRx5ynE2rzDUBsEcmNk/sVS8oTtevSb1P34L6F5
IZ49JIg1F/ENoxd7g+NV/FiWQWypqMFRrpYHn2D1ARLg2h2A1L2f492gdMIlbrw88saQ6dBX06Wv
1gO8+U6QKIaQkwJ3iBvtx49+ac9GUuHFzTHMI7yKSsge5mzn051PJQRr58BBoL+U8yfJFvG9dAi7
Y6LtgYe4eAlA3wIBKdlqCxbpq1OUUZOpFtrOmkaQMCqZZZRikm1w3MyeYAzytrTmkQHqKSiZ/GP/
4IxI7zUBtb/a+gOXX/BxTrKQWKpOz29PlpAbd55O1DagRu+iX+Sv54G4z6s2W9VwjBtapSN+6Nmx
5VSDazIi7eyuCXtXRg5IyCUVFCiv87pIPrqwx8q2N2h+fxM12uLX1x3VvWiGi25ktzaITO1D2s4a
xMg6MeeQ6NncvNq64iKlhiHkRa1rfPUwpTUJ/FtS7IamtdbpK9vGbUyxHf++yI4UKN7NrFk8QxXP
TbHx7ShbPrVPb2xs+TIADdAaJ36IiWuEu9h1xS+JfVS0Ne1yIKigqSxNVKHgibvKqSg+XnlVytcg
HKEAcBBOaSAGQqhNt6hq5y+DfJ2Q2p+T9a2dmDonZmjfeDe6LXknnSf3T1SRG911G3KIZUq00bGX
w4fWp8uglJ7/zgFJXXTQMcrcXhHLWOyCeq4mSAZRoKOGa0M6caThjqXJml5ybSSxbc58o3yuwEJ2
rNkAQyR2u4uFESzz7sAaHVlyx5giHPa2+IEbMa4ZzP6gFNXeWZqi7D1IaHPH89uU8mhGGIZKjVUH
eLi3DT/jrGfZg3en94/LM9Tfs5aCcicBvPPgg6dn3v76zKcRr7Elr4cZOI0fFfuKbRdZwZrTnBSo
6v3ANcm+g/vWULFIl6Qr62q391YKrjUBlDlekhkh140SaQJwf0GYL6azoWwEME+tFVHLcsOhSysp
o4+L+QmZ6AvI3KfF+f0S+h9cIyhaOH63ClzZImbAYtTxFQVJM4/J0JWvtn1MVYETkLtfBpbD72Hu
c/b7Mui/1md8pwaz/wxTnAc44fA5CDpspF91z9s8xDg4x6bhO2n/90WXoSCW9z9ab7pvY2YfWvUa
7M4buMNWdkre7mL54CpOoYVx03pBzGyujEJJq9Cmh1qvsN5OGNVczhbcsVsBpbpBUfOmPved8Qc3
cqjbVYUwkKwi3F8C8p1GcEURi4O1kTe/UsdC1og9HfBsT3nhKVDY0qvL6Ua8d7H2DXUwhu3xt4y9
S96qyBG+M3fehgp0m5fH0OYaLGZEqBkqieOyIrhaDym6CV+Hum1eh0My3Chxhsv8tf2RV7RRaJmd
hKdlRvBntZL+6oxbMtwzbmnqsAWGBkMxTw1JNLwUAMhskQl4QSHoMJ9VfxscY9sdDSAmLYvdxf7i
bvL+oMI7btgfHTq2D9v6cm8DvrpMClbenOMXerZsUbnYjWIgz+kXUXRDKTYfoWGTv3p/p+pSEYDH
BsHALQE3pUuF1hHD/n842c1QJecuWYob4yPMYeukG4dP/iV0MLOu4YnMFY/Kx12FOqTW+KeJFxIb
pwUfnUp5NP5aJDVOxfdjazAcxjAev9Ws3+pPrTTYg7aGWuMqvJHvei+oyjBl98tP0eHXcKcfGRW5
lV70AbHHy+LQO64T664o67duNloxXC3xqS3X7MJKMYRg42fQQT3PpC+mCxdaR/1zT1eCtyB+CI53
qGzU/VIUSe70oMh1mrg19IZcLZzmrh034Gu4HKHZemR/OvY3fk+7Q+kQK8NbfOo0gByXFh6baemk
m1dJGi3BF8J2Ds7NDrOW6Ccl9/2hmVuoVsQOxodGro35SjlFMMAbwLM+c8LcFt7D2Hx3vDw+E6/i
N/mKHBI+AYJ4Fy+REz8z6FjooMlr9PCiaOzgd6kYJ4pzpxeyK74GO6WMdHk1MdgalurQcKFAM5wi
qJwhbJ06AdsqVHoVo9nDyT943a7Ec8VROQho+Jsq1PGjzYuMT9TlmwfdBwyHGkkIxDzDgnMbOZq/
1yKlm/M7R60ltkuUyp8zzoni6YSmcxJArmiL6axmzwAuSdlg6TAPayYb2iA1DiiRSn7/r7haTQSA
BaG7L6ASfjNBEnJ2Ch093u83vLjV/wcjtw4B4CwZS7pvI+1qndeoooqmTD4aWR+3x04YO5I4O2lc
hkI/XkGBzxlSpIV/hR7zRiRXZPsozspLeqn4GaV9Rjs9LLnN3rpHMXEcoCib/ZieBDdl8NbTwuJS
5ZdzavsrziallrUC/4AH5VLbmEyHkI47ajukgQeIu/ui55m7GBpRvyDBMGe7V6ltUJp/BaZlQJL4
ZZURNtF0qYBM/kDHO4fl950uAhrScUyZKAdQdC5rngTw2VJ885VGvSkWXchCRoTMLGZYuOQGCfQ6
mNT56o8K5uFPow26f0YQyEbd0WEmy5v5+XNOo9S4Etztmc5etCVMBwiX5LuEnBLwEzxRkYQfwRkc
1sGEx5tAavecUeliiU0HddUOReeyTJeyy69K75wRI6nws+25QwwslrByZq8UGj98lknxwRkzbatg
q+B/d9Qd6HZPaeS/Fmx41oJ6+h3GGADqJWzlJ437Jq163sazqTtEDaHB0mEpl3yh2AmEq7vt9b2b
0d4buIZSUr9FR/HeFOiABX6jMSOBN3VCI1s8shTTjk8jJdw11TyQ3J7jeb4F5kzXRvN1eh8wc4R+
6AqbalmT09qHjCgPq6p2JNo2dZUWuxdLK6Sm1GPmpRtF7oJJOUDY7NqbG3SY+QdjZrxw5hIf0MJM
5peVrs/etJAtGomVi/HGBtBucgvC585+zc2QEVXCNvedoTrJ2ZGzpyg71Do8vAOyPans26VbD2Nf
ltSdlkY8qNNw6juNwLz0MwT1ayYOt9hb4EzONlSxscSwf9gmhyQdbvyeCN5h1f9XiMOYg4ZO0QgC
O+1/NZL/Aau4KEvzJqN//oYwehgCdjpnG9Pr3F2wgmK96yNm6ia8hl3cat+9sJaAPtRbwy5OG8QZ
p0G1JVre4weL9Pba8M+ShlQ8KK8eaTZrv+lcjOpwRE70o0KqCD9mQtDEMwX/iNSrOkMNBVSefoTg
U9KSzQvh0e41Af34heZvrJkuBY/r0Au17yycbQgeoxC6HTn5Tb7B1HuQI3vT2lHDGTGpMmxL7qX9
q8ss0an7lHvZUKU5Ym7usDY2ObRWYFAHF+pQPKpBYGyhyKKgdS7F0CGLI6ug8n7Bv9Vw6sVhlsnL
AYEb/nlbaANddBnmLofSpqVRoI8bxSEiP+fTLKQlZHtFCXWOru7ZNK7jRVTZEVtM576b7YA5kzAC
odbh67nCSaERQvF0usZKSpE0bIxL2Nr/xFg9ofBLT0570QBbNEwIW6lxTWUIZfDnpOi1FfzfCHtZ
QScmSQUyhsa++GGVOdvqqA+xtpJVgAUANEI2rhAy6UneuU6w/kmZ2g5GNBtLShNgiDIAAs6evfTJ
W8wdO1lkdT1uqPtZ8k11hmsALPd/dUKw81O86qWNJV0zR+Koa/fvGfXgzK/4KIktfiFoJmQAe6GE
WkoyxuW0dlAghcPQzsiln5O+VWdBToh9GlbkRPU9VmNySWvzHSZ5PiRETk6t1fYmdPhPDggzH3zD
ydudPCIlI+Mg4rcUqd9w+EdTLobOYRSvXczbOJFTaPvUX7EcN2VoYSUECpfi/rb4kHec2G19IlaG
E3IM67H9dQd4LmMXzIrloRKDL1GItgPFINzabScf8k0CPV0VkDnYYK8/kYOdgGcUtU0c2LS+CWTJ
hDAjBBzKL5hnyf59d1X59tXOPxT0KRkuodKb4Sak5Tj8B7w3YucY3BSQcPwg7XnNPyzh5y1Kad5M
wV8keappMG2PVcRJhLI05UaZZGwhTc33ZGb1KVmJIWl7V5Zjqh5hwbG+pk+HvJC7RMSzeCpvpDa7
5JEbTAJCFx115bzwnd9JPmUZorQD0edK0v9o0JF43uL+zzUVB6ngmdKpcogzzVC66FaD+bFlEIEQ
hoVqPJKDWe6tl5B3SaY2V69gFr7Tz6OCP9A63/C13Z+nc19y/OQlrkIbXHE8g2uVXZfPQrs0he+l
2Ta3+wSkrynTl1gi04Kd+9m/OOj5Po7bJE63TFYNc0/9Ar5BJxVqqxBzZp83Q6CpcJX83AJ4T+yR
csN5n/InxLZM9wbvtKRWwBI7M5SLZQdrzpFFsxX1tpPeuunPSAn6Ba0Gqv3LusKOm8dzxgFOiudw
TNXupDWOK7GcTrhBEV2L32irN4RCIWurcyU9gIDdG9xBjV/tj8ybnnCuUpLBWAdnF3BYtiyARcHo
zOuC2nkPYSBZlDIzBEi62EkZiLO0XC7uCbcAxC0Bj68XpBi65ihO2FGH8FEi47wb+D7qSUsz0bxg
94CcfQX2iRr/sTfMzEnkWWPruSGZNQfcc8H4QKmuclHi+yqOqKg4rXYF+DGLVzqbtp3Rowr642U5
9oFJmYBtpFcyAtgDRTM0+riKtLJ2ILLrGY8U7jpSuxtO8V/tjSOrK394IVLlEtveVwlzKIS7q225
zNQ9/h2VmIYVE5JVc45q9cVTUqeYfvAn8Zfb5epABBzDHtKryrEBBKypcNB+zhlQTKEnBKulv+ZO
Bm1bRbEntd6KNVVlS1LB2WZ646Ndc2+asW2axpDGfK+SSAWYfCmGWXbbaB5WQj5dORjFPMooX53X
/X2NwPK5f6Q+NIfMSOzilyIOu8EGTm80FnbAGxHTCYlTa8amI78tbOnWD1lFCRAZUP8XdqeyBXg5
aEu8KtcVfE8GeWMYtjvDVgODlQWLghhOZovbYWYhmVCJUgOwAXdCJB13CaBF+V/4Sibrue18pDCd
20rsrU7HAmysAG7M7TgAyEMl90CHKxuIzfE7inT26YutbjHPIqyK2wIMNVtHyXbllqMUUpApRaF6
7ZIK1PzhKLAhE+InGHeqlK9RWEjtlN8BFEgJsKI0smqinWOEWHHFYYXUQ7H/FdMN6SYi2XCpm+Xl
LTHgZBfmv2NwqQrf39TyNCbrtIoYSudS4awXtdjF34TXKKKAwvLf4bIQIPpW2DsA9s1Qupj1KORs
FKJwLmSg+A99/izklY+50m/IWtLyEjKzTrDYWItsXGPhukjgdqREOPEBzGJa0hLKPBmhJAgvAfvH
qsJ4EzRL3VQvogdIOavOdpqVU4swfuLQ2tx1x4Rb6Mp76RCz+4on6IphnQ8qKy8JudCKXYQbp9Zb
gpxUqNKln3OlgcHIZgkx2liRPmAUnVZr85u79G9tMoxmXyX/2SnazPBiyDlZjRlxciC/vsj9QPXU
o5pPa0rCDYPh8hck/hVkYJUZiBm/se4d8hdA80wozKeOPaOSRy9bRyhqooF4vGyP6h8n0voOnSPG
wgrhiLUfF2PwBMRn4obaDdSoiMio61c2bQlkiPV7owiimdeWlMVilSgDIiYaV3AuTG6Bl0Vnmphb
Se9oVo4qPJPZUIR9hWVttdb9Rthhkc1MyvYQiANRL2kD091VNKV1z3vFtcZTFILV705EykHLBefp
kS0TS/0y7zkgxowLw3wAwG7Z2W2r+YhGEUM4nLBe68ak8gMsaFEMhsKDnet1YKu/qHeWdg22KcYl
r1S+x4uzNTV5zU3Hl5nASCdW8r1IU6HpqAmHZn2603n0V9WlQf292cMR/EQY9JTdogzGrmTALA3Y
4rt2ipymCUuqyu3k3mp5bQ+f6q4qzWDCiuUd7VRBRA5iGldsqIxyoOEyyuBLC+5mCjxBjkf/O43u
fm1M6EtkH29anOlrDTd45u+HskbcAJ/7pJkfj8fC5XQu9eFFbe3qRTaGv5F5mVIwq2y8DXrIPRGf
iCIyDtSLAJEuD6BJt3WoLgR8ElLPILItVsXKQCRS6JjqJuU6/qXu3tdTRYeR6unxXboYYsY9v9Vs
uPOOnUGrnEalt/K/kdYnunQjw0+vIxxSFUghLXhn/yOKVwbYY359xLWJq4Rn/w6AzxRRd7vJmGq7
gZvnwA9jOPFWTWvDuhQQmCQh3tOui0hGqQP1HDsLa+IyJKkVjXopS2kzTi+ge7qNcEbZbW5LMoLE
TMGTcxJmMmIcA1qOMf6MLLWNcuqp9DsSW7Bm+rJVD1dE9niwGEO2+1InzXtwIdScEayrTaiSLNEZ
hGzmYkdbbeYVH9+Ulpkl6XowZP9k6rA9xAEOdvSmoNnQVDUm6nxg3q5T5gvaRiC0ECrrc2614ceR
gKKYTUDwTFCYzhNMNZpTuwYaE4sBPEaWcFf4vvbQ8UqyM22p4Ix8ALTdGkNcH94Knjw9ZcnCZrVu
RNp5whBQdIGqNKPNg3PiiN2SXfsQm5u5q903/FGJIsAOi2sn5xHemipW3i3KwRbhqaFbyNscPivv
sk2TmKVvq1Tz+O5AHeT3MxBfO8MDmjw5sXlWi+xSSsLD/FcYsf8IcNqIxX5Qx+/241hYbUZxAL9f
nZo3lEplO68Mmtv4MES2APBA7f7G/zD/DTxj8iSCDqqFZgDEC6a4k9FntGifHFwZ8OhgPmbmI0IR
Liq9ro8QrPJXwIyaGfs7iewU6fu67mRSzEaWOi6W44dK/fEiHKQA6RhOx7FXKKt6WizW7Yp7SbeE
AI5av6FGr8jg1Wlu7rXyt/k3rZh0Xu2W9xxlnJJcWisRE5t/qCmSctKemLpLMBOfQoQg9/F/Gbsj
cXI2vg6mCLb2p1eo+XBNRyxaHsmbdRLmVxcqLoChlhrZzzyzWvWIYZDRM9IRGv8iXd6F4nzAzROi
S8ctlHAhKvsz7SH7EI3fm+JEJcUl7KKCpe2tww3W0v/9ultuDquMbVfwL3SxwL9AXAxA2bQhY3Cl
aDiWSWzncRe7c2OP7jhQqISVlK9ho1cfCLwOOrSRCf7JoUEoP+2EqV4Wy5NoEI/qQo/CqKE3rh19
Wj1OVNOiiY4s3+lDRtut0bseU+5rn3W6NwycnP0vS2bbODV+ZQ+8PtQgX5jkPx0NJspUw78DNsPJ
LiJawkMtFeKfL9p+wzQCVE6NjzvdYNp4aTu9/hhs4vNKYIjdxz0pfyutD1tAgnlY0b1/og+QyNha
4lmVCEYV8YjK7RctglsLz4ZiG7Dnn8d2LkaM7/3dRWcCXh0GU69es0i5UDnu0LUryGjFIjaKjn9w
uiFCE5r+qRFoELXcDzVI8XU9W0aQVLjIhs9DtamR6kkQm6TwNMZ3ZowCgAou1C+Cr02yHWDfwx4H
l1EXGmiqTjeoo6LnJpUNWVz5lOy4yUWOe2DPYovwwJDixXS4wb8pb/rYfVcblWh3nrNi5RKTv7yw
orgCVqc9lSef4X+/JTvWWCJlGACPn1RCvVwBg56Ch3ccwcucYif8v8sQ9/8Xjooc9OSVAFMOs0m6
fbSYbi7wz8NfegvvAmD3j3AY662w69bu1h6xPNPRjuehPhHTygLbr2xui3c+3F95kFc7mRQHm460
M+FFzh6wVjEoTbMIoHiCEVgd3znTCTTVcDJcUqH1FZgAXikIxtV4tR24nQglEiW/H4AgeDTw9ALc
R3YPiX4+Tyttja21Yj+vkTrXt34ZJQRflQRjvGiEYANk8Ww0AvCnborhUVWh8yiFMsNyla18r6tM
izgwPnoQbrngGmglW7yhrfq5Jz/JgX8r4xweO/KD48HGHTryWJWXeT6Q/ZogbhidlkE2MeP/Lh5s
byR8ImUOhvncdxvA+CcqvV7oujUMAOIxYow52uvp9zyQFjKNju3Ls3lbCFiib4pmKWbE5A6d+rXU
LogURWTOl1R1UekI/njAm4+htb7wp5LbX7jpFtzfyrCVI32w20L4a5oRoz8STGPsACHYBcq1jK2W
2urIlPnAUUMO3fss0ZeZQO2CoLL22ozhqpqIER/Y04jeWWleBDGfjhBYzzSa4MQrjiYUEalZkeSd
2b+OzGxscIonDw7wIkTndsiQE/Ad/h46D8vQn8ppWqIeYeM9BoAIQk6EVa/ZSNMdfNDHr2UTfnOV
KHaB0FJstoGj6tipzl8wa/sa12TQHGPhHXwWBVXGIWy/ADLUFMGwoloygErrpRXrODGWXV44Vusp
f2XxzJCjcAbf5hL1TNczT9eEmh5cXxnbDH5WFDHTsC3iQF9Vrg3fbiW0tJRnvqSD38Mc2zxJCd8I
nPuJUuZYK03VUVLJ8sbIBx8Gbc+EVzgXt/O1+znJYr7u+5yF9ZydM2Bk5RB1v6uiUDXN2cQsEJx1
KZWeGBUn05Tmf1KsoiIqEkjvQSZv8KSECyoTu5xsfAbaiqX37oCYm5HsuTTNIPGLvTooNrUjV+LN
6qxCwiFF3qCKXVNQxTxYDkL58jqBf71EGEsAq4rwXqBNb4IlSAjoNVIMnW5tiDSRJOus3f6MLzY3
rBwcpf0b+56Lw8qb3cHdVBxXj7WCs0LFP/jjr7a2Sb/T32OmZV622lI9aDDtWVJdMcK24Lv5EMeT
4ZabEerQwIZPhr1DHaF5xj/wL/S3QYFS0xo5u6CnIH+uyTDBEj6Q99DZu+m3tmNUJjKva0Z05Nbv
fX0M0TloWo5e7zdcKN+fSCKJWuoYGqE1je/AxUx+VX4Dm7Yqrgw/X/54JOHI1A7V1IOFqUj52jgo
78WWHyRbxWkdlitAGPEfRmaH09/AttDueHHPw5NKjqTkayl0uwdipKa/iNOrwq54jSDPBPBQ9gc6
2hr2iD3tvh9MTfr7HgMA+F8xEH/dge3oOdYUCfgYv9SOWl03pgWetQPSjAQUIUhgqSnm+0nHo6zw
1SPEj/MKMJLEoGU0d0BSJWcR+TsueqMI1F/pRh+ND0PikSnDm/2gB+vZ64dNhOe/OvL4y8juMdR+
IJNln2z5e+ZJzKqgxoZcWhRg4f39Il7a7ArIIrCECfhaO4YdxHQqBtIFRvE7zhAQDLhNzdafqYva
wChxfwnCQ0ZNlC/ehMAssHiv1GE48zxqBWdO9DxqSSbxrJsoLYQACR0sBVToQCIONnz74DoGORsa
2/UXBlOeurQ0DFElYE/6axQpoR2zcajOstVUmNLvJxD1ORgZEfATEAbHETEmNI/5QAP+TRySHCAa
ZKI4y+OiovjXtcZtxZlaej2yRQk38+MCdL93W+GOVYzKpLAbrspuMcrII/EM7oGwbSMToAVKt9Qv
ORHVyWGSzBfcLt6utHjuShW3RocPBm32j7uKBLezmaLeYAWj/TZ16VMLTr8UiQCC1L/gKNcOO+Vs
k0mkfeOh793EQdetcRfqkv7lmc0jHLkZ6nFz3MTtnQAZEZYtRYL4ZxZVkBYba5lhQv0cUwodbhal
CfE0DTelTHZbWsdlAj4lpBoZsUanP/A+iPhV+QpXqk4c10V45eQh4TFSCa+/RdMLdXt7B9K9WbQl
yTIYL7IvOAtF8bSmXWrWOzrzidmduLQCQYhCxzzUxbof1PFkHWPEYTj1KSyN80DpTfklaEVBaJ54
gEi2Eq/RgjLzn36WYG4FBCudWRdlpQLCCNKv+U+Q4m9O+HEMc4/K9HXrgaMwMZ667t5KN6aVOpJY
aGvvKLTNeIFAB4+UaTIwdAwZItuCbo9tsNdw+pQd9+lmcXFHFO5xtp4J39DSg/JQpL8a2UfhledZ
aD8I/3gki6sU7QePyKDq0+llRc5jggf0pHfGrs9kWAe41HroZLpAb6fZMOo4Zk08IlN0engEKk2c
7UMUO7l6U7qMtCOWtmOdgz92wXgRNa+MRTm3+oAD3C27xgdE+a6tStgzXfpX1jOoZ4CltUwq9jRh
RItXXRgXw8LNckYMTDMSqWhHa6c5s5Mw60WtdsC5PFy3hnEj3axU4LYwMN7uIkCc9dOgzKXrGF/O
MrUGPQceNJ8Qjm4e3lNEgirhPLeYPolSXJbjxxAUwZVr4cy4uoYJT+bYnqJp+T5DXIgwS3vvWIHQ
ir0AgwAP+FDz+6jb82CInhL7rMPigsz2CwS80P03OcD0l7YyZ5kCFj6HTHVv0C3N6m9Aj1mFczX7
2Ej8MmQg4qxl6GNaO3kpBgCjhSvKse4nbKIZbmSD2sIrRfl5/bDl20JdOUpB3Mfi7yKluJRcLrrd
mXOi7pp5P/0DnJ4D4Tg0e5XkVl0IZ73cxANxfFTt09exVmOPI/BQycsrpT4cmJbZCaMyy9EhlJT5
S9r42ZpUM8nbxchc1acoROC4dsRvIQ2Dd4wLV+B2oKBPfCE1/lXDaWpMGPhvbthZN+43iMt1RSVv
bRp5fqg5vAOaIUUZC3eKL/9VWcdRZYI8EG2juGZFt6GWYJIMiHyr5QmrbdFjsvuXXTO79hHaejS0
g1aL7sdgyHXslvlPHKm+Qh2skH8NK9ibsfgpjF2iYeen3guPbEBhujy32txAmjPyVEnzmj/pjMyz
//UV9Jd7RVVtlcND7oDdhFpoX3tkza5NFMZdjSwuhmFH7KnSB+c6JHDZTLc+6HAGKj7/ND8FKJ3T
f/LhG6LC6IOKwuKX8gTjferFQcHbwQ/0jn0G3RJSeG6TYoNTq7lCFgbMgX9o0l1oUGWgoI4WZgQU
D/j/w+su9ZcxCEu7f0vpRlHEDK1wQIyFNq+7asCOoxTR79j9/gpXMFxFWvgbUb78RSnjq02jCeFn
W7xNy/J5LC757fc1+w9svDW+xj6TcYi7KFWH+3gmb0pPIg7tFwGq6N5hcXsgOkPMzHpBFIcwELP5
7O6vaBBrGUGtnr9UoFOAmufKo7q8oXHGFVGI15OTG4rWVygB3Zu3GwVkM24AJ9/L1hH0bc0LxBY5
lp9t95k1WZOvDTB9xjyu2wHgesJX0TgoOeLWob/eA70PQfhf5ZG9vuJCjniYORTLaW556JGsImP7
eGM+Hn2cDFB1cIKmDHmssKprK/XXODuJuQWdo9LGwwjswzaflsn+R2YR6ej4Q82DMHJYaSZH0bim
pYk9oGD8Wk2phgXA7JmRmcmZBfOrBWRBsEBxxj1cQxASD/5yW40HEUCPhYvmHFdrSvgbldPAVCvm
suJUNlPsmqUW8vZER63ogfCSOtrmxyhpvZr2ITpO8Q+UvYBVh1UgJB5KksDDro99NOHXYexLbZzc
uqt42/IUA4uQ17x2ZvfDBcbLYXYRcTiuAsm+i+GxZKsdHXrn+M9OgRZj6uzs0wC2IkJB1aEDySgv
+bN8GzT/f0kDS5j6CW1n9h0D3k7ZnbA8FAdgiGCzAgLLjj7P4W2M5SBQaDiziH3TaQgk/4/3tL6H
vyzXzJT5ICJAbmaYYo5bKGPl7wISR5wXkH9OpzFCej8AfvieMwnyGv2DcPOeE9eZ7ZfMNbW16sxg
eIHY7Xm3POACpnweIDPMKsVYM7X0ULy7eC4uURr2Q0Psm+2zM2x3fOgGQ1He2VlyHHwupxxVHT5B
Qf0npV/aQa2v6iYtz+ChKyrg5dFnshOCj6M3t+uhjR1zejBUrqaSsseIyEkd/7Q0RhYBRrPaIe/B
VVTgNXnrEZenwajVhzIcuPTv1UQ6bMwxK2EX0RBkY2+9030fxJRoniVfdt1pV+DrawvGGHG8ndQl
SX67yO0KohhXwGgkigT+++15TMpJC6DT+F/+NZQAlDxGC0R3thRwLH47nlJvJcLXzOKvDyoNVboP
IIj3rQ6/uxlsuPh9DNTh37Iid8Rk8j54oNgUMAhARsGTM0HVZ2YsHiSapBD8/ptF70BIps/Ps0+w
AFf1BamBjnromg+Dgr0v8wUJYKxOCDcQsh34eZH8CRAWppa20Qyvsux2FPA4KJaUSWiNn3DFycHm
RqsDOrjg9FNf++PixUwqHdGAUMdKPnWnl96G1eiOVq/3jOiDXMPuD0ols8TYiI4DHX0bHHmZ9yCT
PfRq5GTAxPKYDNB3JETBzlYNvSKI35Imz73044JqhoqGsIS9w9WU7/hwN0QMYdyir1LRYf35zsDr
sLGzHPi6YENImXlW47WASj5iurdLeBv5Hua1xyWD6V9uf129V3SMuz6a/IpolymAlrOxDpi45I3p
jtbS+JAaN9RvAWOGT2NyXmBWiERi5Zy80RYUbjXBy1x3PvFIARGPzUWTUL0IrVX0+N+Wb9da7kCY
lyN/EFBD0k3iE1CyV8jKJVanJNnHtAc3GkgujK1WXoHlcuYN1x3KpkEZLORQkqoxMNVxB1cSNJbq
3YLA8bMVGzyI4OiWAjwuXp1l2ygJZXbYjqFPGR3GTd4f2yEPEIwbMXGFSbRTTDDgs2m28kqb32TI
AEAYUIZbHPeE5dDmAHK/L3TyAY6ORNkKgOkKo6+YLRp+xkYBJjSiAJycUxe17AffROTOiDw5t0sz
j0hYHqF9QmdFzeqNbNGdizZd3xVOXExkTe/EWT+XN74S/KEtKb+tQv27tAmNbIaDhLGnpBiHx1VY
Ooed0MJMeM/QXj4BtOlDY8YsYAp+MiuO2Wo+OoO0/M+OQS01NX4i6Dm/I1cE3sFiFiMSfrpCzzbF
1Nk1xxd4Ny/UMcxfl01xxHRVrZaXZOCramhaccRTPDvfr2hgkYkR9BZG93eAURvec20dQk9PWiOH
r6vV2f4IDBwsADWFG+w1oCHeZBVPZJp/mobdXdtmLDqanJTPWwqozZU2hCYFq+pl4ye7X9MZXONA
/KcVTd8MJc21oKqrhSdjJz/VNsKdGXG/wcMCafYF2iRR5TRFW6lYA94jrKLEYX2jwnbQVrRfZOGK
d0xrqahpecyjJ9hFAkBxfWGDQ+MWGucDhGas9SY6Q9oDFoGQImIujwQMVo0SC2UWFmXfR9CapzJZ
DUZ7rIuBpBeLvM+bi8wRzGTAO88hWi3R7Fn1LdhSrvzjHalBj06NiACl0SZ+DOkc+96FNtV63QMD
ErfuqHCmfmw+ydwQV2gkVodBXjVmoMP+k4utXL0pCQTOgAkRcDQVcBjgr8H3X1bqcO+mj8gvnPfL
Bq7lks0eibQPx5QjVaDcON+o5xEz8bYtmJYkWL5qhXVNYHWSYeOt3wFSY6B7VV8+Z2PLGKkqwF1C
OCrqAzPTDNcJkhO6DEYXBWJOJrwtISFohvdhn4euEGx8PK1Ai2lT2UX6tzUmfrwR9k+fz/kBuSCB
WJBYfZW1p3upWFpNJuDOwhdUJplglqQCkqG4S3lhIc6c0WUDvZXQJlIU2vgHgZUowtTQVdmIqCx6
6g6NVTqGP0WqZkoTg5gnARqMCkW3ML2/yXCUZEQCzMsbw+PNrkk+higIBB2lVIuDoZwSwBuhrnG6
NVTJk8AXncEllVHswq6uMJF60VGTN7pd4TT88hGljhlfmZJ7/hKcPi8Io+Z9EkaJ8yxlDDoeCzEr
v8pTqRF8asrs15jaTFixSKkc19UB7u0JETNyM9N4q0BH4Vt6Mw8Tzm6TfiGDOSnN8KO+WBB7dyfZ
GdclBa4RdIOGp6F7LjaKPMM9QDfjbgD3U9jjblxfqwm5jyb40talGcUK4gtKQZO0FzcF3b9ojhSM
YGFgdZfu9JYW2YL4UwBbIiqktAXSMv2otwqTJh4dSIQiQ/u143GC8cYZRBX6wRGiGDlfHQzbeoJT
AglxiJcrw9kGMFKLoKwWQhbLSZ5ewwcfti7ShzCJTLGefwzSMS+BrdjMuDcUgPHQOBhCe1oBZcZh
bEINffKz1CLUKpmBgrQYNAyP+FKxnOxAwnFxyMEYK6SY1ouqXhR0dyC/ObIILP4x9JQkKIc+2dfP
g4qB4XU+H7e9joE4JxkDRgjODiEZ3aC+JkHMG9itkdMjP2nG1rbeXRMgMNy3e3UJS6iqF1AEQIyI
Hswe4nctrIiibS2wbEJ1HQM7SOSa80PdbHAdulFCuw4+dltLj6qobb+e6QbLv8E7lNClEWVAIMEk
eouyLXjY6q1wIEh7rLkQ4R6+UQUfLkoxvanzRqplG1zBGH3YfBXhRdejOieI53RqvGIYhn1+qvbD
8F3HRufgDBQ/yiGkGzMgQoh+jnf5tzTTksApNINYOxY19jkSI82ZrNaakryK0YvJrGwjHqDZnerb
muMwufiykheuN3hiVKYdoZeNtfRmW/9Nf4bruIAiZ2pf+Yk9MU/XbCRjYgfSCH5ETtfBI5TQQR2i
FoioBeeU+cIVIdaOGNIcvMspi/RkA0ekBp62FqxVjuhbDXXD9S51p7gkk4WtdgLmqCgJ6eVXhBKG
TKB0QyWnYCQsWKFOerE4AlLSwfaBa9SAq1F2JmIik5lcQh8QfifYRdH8Y7ZWxgUVmsZUqjp8UzJS
FMfYDrG9uGplZp30QhLBzTEDLjHeRddpFcJ9oMK8S9aYbXlAqAY2YKKUQtVeQuxYecb6X1gg1nI3
vCT0IG+0oz80AlKrOJSFMflaNBjIEVn7yW8Lv9UcOcHmiWRb5kWAXCxfFK449wY6VZogEUzF3i9g
JTpkvJi7cLlREdkpmWTrQ3rm6z2OZ/h1wdIGzPXL2qkJ1u99ClrRbeVBKhl9tRCBcOKRbMejcgg0
M2E2cS9+WfwDYc56ExShH5YZA6hhHpxF9koqErJpn5Z7sdkqcNy5XMzgUUYYMUSC3e8d+Wdepi7g
jrHg4Sn9MAjWSgdm8eRfgFC3ivK79C7JbPbRewkQD1vrdlf1ct/7hvrf2XttIRCbRwuIOCn4h4NV
3KD/M/DkpBaahWBFBbuaprobf0Hf94nFhp3ERDt1mpYZthN6JIqyCvD+r+jTBT4v6jDveOAkHQ1c
4oho8PIyR9I3TGsMC2zTZWZ6l+3ZSBzqySRxzl3GHE/deA94RnRltWBYI2rgXN/wSjVzVIQxUtr8
jW+HFBufCFakCaL6mUAmsg92i/fb6x+BjmI7ctzB2y+m40rGwa+7HiITzt1umpX5NEAji24BPMNI
MNgfzjNNgFVUfIOMokI7z1A4182pYob9hhPL28eCZmhWonEE/5zUVEDFIhmEjF0cl0ACv1XY37S+
M4jrHMHgzU5bAOzBplX/PhfVrRRaAUCJU5qnzCGql3yDEfFo6STyoVS/6Cr5mE0FHj9aP96Y7MXN
hXS7JXxDS9b0/7JFiPUOnW3Ngu/s00kDLiboTpqSGVKyxq8WskICWCcDM4arr0lOSX+wGv2etm+C
gmRxyssaF5qsCh5PfMWSN43tjhc4FDBl6YnXmS/Q8Yy+ooI5d4WM+QyCUDwZW2mjnJVVe3VncJEo
xtpvshtM1oGrV8goMxAYPevyOiOoHg/seOf0KH+XaPjNZjUuRnWFcM1n7vN7cvfS6O2lbiO6EXpg
BW/wVlNwtvJGIUNWA14/7JBfexf2/nkca5bBHOTESB7Xrk2Qkq9dieF3al4qzGsOl8Aq5iMpFi+Z
56tQT/jfciK1kEXiNoX9Nwpl4PTe9ZFaMOQHnRBz58aJceaXUd3QISL6/R5AMYEUrh3rMgWXaNjA
vxx52HkVdUufWY1n4EhKUylekQ2zB7irrxyyuS9lAU2ArHHP4NzRsZT2WMYOO1Yc6QHhsdLzIhaR
JldI4xrHUoj7M8dREEF5NmbUwvxdbaG8Hz1PAfcqXYCjHvDvejNVOdohge4RoqO5PA5K/a9mrwR/
lUglOOqbL7pij4VkJoJLcqtIJhrKyhipfsi43mBhbxWUVbivI7nr7sUqoZ+ONcr5p2QWB2OTVwGV
1Pp29fD002BK/HP7q9KJX2oB6ZPEeSmKVw8JED4s/L+7HEjh77VeEPTN9ZW+j08ifk+a2obXgNAl
jTLPHNCPXAjd0uD9QdPIOuqllGKb8eAX8ag0ggBkDBye6FmNGk2EvNjoBRADuSL6K0f8/Rm8lyVD
r+tjuyoVAfVzEpHcTyX8N6Sq7t3/wdXjVAfHgKrKsFWDJTCxJZWodls307eMiY74Ebjg/hcG1hsJ
6IQfPksH7oIEu6XOb++w7irpQm5zI+VeyoKxVvubsG/KiekYop750qLxqiAkKndxNv6Opb4ETDEO
Rv9WEjEfyyC7KKhU+lr3Jv+6ml9G15qdWSXq5hXO1JH1St9/HM1EY1GAbrPVeM5m2k/IPkYVJghD
Il9Q++5ktbNVtYl2IkT+g7JyzAWN96eLAminzfO6v1xW5bFsA/xW2tUgdH+hf584uQyjtPJ6aKQA
MGuNf+FhxOOX/ZIJsfIfbhQI1mGq2pmmH8z4+VXCdSdEWcIhm9iy/WkTic4wks19X8lR7pPbJbGo
LBT7Hlxy60iktKRGYLjRmgMt3z0cJqqncMYR/K8jsVTpITyB4eAVWQZpkVFq4RMaXy+rN98GrOPG
X8vd/CrQFPUWIDnO7s7YaoaaTPvvp4HLzqDacPCxUKhYnVReuw3U4I3WhTqYSDG0yEJpkbe+g5nM
ZqQIra7bx5moliJ+mgDF/Tej0xXZjBPkooHyGeDGH1SVadQHIIBDl3OtNtDTVbhNxeyYpwdGS4zQ
6C8UdFRoc6UQT0NA6fc2QYc72C3J2K9lcFJUFnqyhZ3KldBwOUQs2QbsioMWkVzT5S04PChP05jn
0mE+obmjCEzY9nSBzH8x4tCxbaUhXmF7FOS/+t414WNUZqxy2d94EayV6FLAQkLVIdA7eHjOaS4X
FcfGtqA6dJUGiJQ4/XEmJJr4rrRarLHyVVUNPERrnl2HCvWpxczTPkkyZ8JpYy4FsPCTKFxZyXos
xitMNlp+DalKpVxUpgcU6m997veX3tcYqUdO9YYTI6PR+5hYOCHXijvM2Nhb8eT0+imnAQQyc5kc
hdWxXZ3YjovICwH0T474x67lxuafVSzimInYkReXmHpVpXkFGsmfC3Vn+IjeyduWzhC2frdMHSvq
AwS3HoVxbZ9iG61rqI6xcnbeHewGjRhazrFAi+dRHKr0c4qBb9PP3zZLyH+a9VMEiZPjK9vfOmjQ
H+YyxtYdW42N/cK6rSSjK+vBH7tKrIPqT2GJw2ZqvFCLY7rfq8/SZL/TIk+KLDuF4FShzBTUNVOf
vDThhNorKQMh/zq2NshqwFL4A90ebi0zu2qAkVAVY9IXj0hoZw6bXOVVSoGDJR6KihiZWci8dtIs
EkqXdL5Ybk0UnMvMppRk4kXS9HBgDsPjySHuTFdX4vMNuL2WrqeaiZ7U1qOj92VEkKX2dvxR7TCP
lhRE5mqhlpB2EY9Inuto1X4X9Xkz51Zzz7IP3aWxDV9opayJeDI0coDezc/fed3UxLaW8qcuf8v0
YHpmHqK56quFOhP9b8xzbH39A9fuSFRJ7crtLc/e/DyNSsusSMAnnWwcY3/MqkqXJVQxp62sQZDn
mkptjo6bsUFM/nwBOUcVUmwzcd/w1UY/Vr4VFbwTirq4blQum58v6MbIF0JnrvnwxQUH1+Dsa2mx
76BU4FDA3eAePIhkV+luMUHUpt2kTcxm/AN4GKC7OSdezNnm+iyCkARQH4rXtB7k3yMrdf/YOs5n
k8Fv3CQ5gkKKXoy0gDhhncRuWFA/OKpBsRxxbr7JZJpUBf0VvCSPdatywUwrp5htQCVt4gLnJt2x
nrJGxwgJ/oxQG7kHPpE1tXoVn48H2gZ2pJVt+zyNJMPV4jtSWnOGL97er7s8vZANpfAIWXHNp+b1
k9o0mLZyCdwLbubBDgV9qGKiIlwkXbXNx5rrwYHBOA054sJUzrbUDDajnYGSd0/6h65mSO/IdtUb
CPEH9u88o8M65T8RfBYSoFRBBIdR5m55UFP/C7L35AOCANtDEI7FMYHF9R1Te76oEWrK/H8LVvVp
VoA6x0S5bPGcxueWJQ+CQLzoWRz1cyKEramGbn7ycYakP8QziSjJQLtsVPXBh1ht7wU+PRJL5HWu
0I2ezdsa7d2fznOnsiqkcAfpW7eBY0Ry5hzqvBmpYokrriGIAu4g4khE7YQ9o1MhR08zlIkmhlLe
FcuxxaV4h6Ty1MQcKtahhz2mJwlz+Ik0vtrwlBpc9IOcDF7bnORcQQ8ZqU0I3nBynKpXjZpvw5Iq
6md6DZ/2vUhHN/3RcqPjWpVpHMdP9ya6JOQXxuRIVYb/MfYVGz3d8EXNxNXJfBpipsGCfjsKMoch
oDD2jp4KEROVG8qq9H6bTL5tWdqVkBo9pDXKHyzBGvikpEKGHtAeJ/L4DrWOqeIl3w4CO8+7ki8v
T5kH+dj0GHbk1+j9V4TiFoBLqmkIw/J1f3NoV+2tNPBt4tN87I7NubL7yf4avwif1sGr374EkjQL
pHwmfTrrCZyhNag349kNHz1ZDbsm1sjvSvPLj2bUk8k6DeVzRgakFQmYbZ+iZMHgdhZX55KK2A0A
Z1QGdaCxyYLyIU53fQArgmbAaoifpshJ67+ddYENK5DFO+5+dIOTgFq7XqUjkPOZnf10HHU8BSxZ
BKYolX84HGmzHpxKgG18AqISqfnhzNFulqeUCTYOGzJpdkWwXSH9J1Jtk4AXSrG1l3MshSumc3BC
ttpogss9BPs9X2pmDaE80/7HTxk49hZZPUF/Im9dq6Y3tUmDQn2qB+n1zzxP+/MCGpMZ+l+6WnPY
+1DvRhyY3ejSlrrqlTSy57Cr7wK5QDnKO/IG5XUCtzAFQX47zBsy4qOwXyiJsx5pUUfLQVLQWuqJ
iM9UwqlkzZ11RxU4RuzpStg4TUD/epRFEvZVHCF96rgKh9X0KqC/5nZsPEl8dzWZa2PdMtGs48Zl
qXkDrh4OFzzF40RzP6pyKC14SqpQDQL5oB+928AgUSTnEtWCZzzY5q+vHccBDKz4QcRamAiTOJmS
B19DV0mwHu36512ncpnedBerXgDrChbJD8DmWOe+ERNtnvLf+Awi7ct17rRXedW+tUcGDIrK7U25
lri8t7ri6CyE3S/w4fw3dbq//Yn36byqO2qLHvurHdg3PEIJx+xICvXgtCz86/d6ObgYtScInKEI
4Vs5vQp5cornPInNgAlkLmk61Y8tsSYp/SipCeYc53ha3ZibyB6zaltDnjyhL63Kgwz70vLFavWL
6FlV/0Vv1E6iNm7ZkgyPBHyMx65bzhVLHNXHOO8QJu+Q94ureXRjPD35mTe3Jg4QkUTmhwwNwGI0
HnjMP8ksvnRM0GT2lM/M4VeEYAlWNaE2517aHKqKOYO6lIBY7tHW3/bCPpEGjmwBpNMoNn4WCi1d
ZX6xjCqbv/xoi7q+OTJiWWqvk/zpJ/+5guFzLaP2k0FU4xcwiTKr8fHPodKUo+LHO2Ss/Hpe+uWO
3Ro2Z+nUvwAF34CdTCuMqU3+U65soArcZAO/BE+RzQOVis69Ef07j2C8tgGzcsJhpHp1FwqO5TwF
kc3auJd9OSGBdWFN2RUgKIKO3wQ4DPCYsY2eZ4c2XzhV3Wgk1J7Dl8btweN+jpO6ehyU+VwtraES
cfDQ3MN7kzQOPU9YMe4H8T9PP++82DjGOlmv+YpKq5tMcu0dlTMOnrq4KESFqe3dp+11ZndFs2cD
TRut28F7McorwTG7TQuy9Q5TQZLPPK5vU5loJhtfCNuGJrelQy7c7e0g3RSSE2lHH7E0/+QV8+uK
JDZuxRZBC1RXtYcBUk3N3bXhbpmI/3y5p8V3m+6w3iOMAiiHqFRsf+2xoLctI2FwUkxDkDVbgv5F
2/Hj1PcisUJ00g8fTkH5ZKoPjIUvtS4PtD1wlIEwNaq5vTK578NIKwEeBiCCG7o/wIxhveBI3bxr
8PLI80Y1+UWd5WhwYf2UciWwjaPU7OSyRqOspS1nQDkVPfXPLV0fiKRBiuNcp3dgkzHP82TA4wHQ
FUSi/27iSuXBNk6k4wfFFFQbBW0BnsKXCq4mzNtA1WOcabUMwfqDuocuNqLVw35y86kX47PFat3I
LEIoYi93r2gxjUDon/l+YZWyTo4Hm5Epc9rcJHcn5ymFgcthEZbVZs9WAPlM5PIAvcbUSlsMzf1V
m6qbvntWqC4TW6VuAA8uVILAGaUOG5xDaF8kRGQr7ZnpZ7KrE6ZkfGZc50Jf5POCpXOELbJCcWT8
CaFtuvlF9G2349/1fE0ax8keAh+4iEdN3Y5AAzCzxCSUmPXnuY4vurNA+JDmVLHxrHTFhm/yrAPt
yxttMQ34NYwddG6vUUPuoR3coCr69TEw1lnMMhfxprG6M88vnwjjE7vrFb/pynQ86Nzo4RARKlmA
+7jOt/YpmL09MEW/2WTwghHhkZqSmo5mlsBVakrrKgP8zyv4UcaxKaobSmN6Humtf5XlAlf6SXIu
ibrsx+kKkFd7M1iSA/hqHU960kwpTbwxbHwTHzi2fC5NZp2XxiJMM7wE2QqC8Wg7Jh6pL9dAEvjF
4grDkXIO6TfUFdnntP0A01D1p8gUZD1oYJgXyvGJU1jtBlhOjSlInTeonik0W9DCRSTAKg87qtg4
g1r9MLZXgYbboQt/axvdQGhsiD8AccU4zHQ2u+wpnVhropEpB9UP1mV3KTwQJnYoPOpJZWgySQ2+
jeXCKsASHsl9o/ZiBxyVPjP5KVIREzzBK8nNhgj+W8Uvb0AGM278r4j/CGgzYQPIRL/p3KNTzl6T
6KBhtOR4rwVER/g6xXTQYxCeeAy3BldcqEfXS8outIQ+23lskzmfnzFdEu6dZWBNCdx0hOKyFOzs
cv60lxZ0lnLYV8bVLTtCqTBg3+AOheuZs+ewjbN1GkJolxW7kepWKCx5/82sDxTBtu1LEeFL2teC
elpj3vbcYWwZ96SXct6Mv0CZ9ev+uMgWmwKcmp3NMQmSruRCHMIaZSbt4Oj97mpDEUBYdyDHMr1E
GeA+AKW9i5D18/Gdh/cG1ch+K6JOTa9muXyB0FXpX7aUjdu8O9MvByLhfROaApz5KKVx6Hwogjzw
Vl7cGYX5bPNa3lNKQg4OOjMKBeq4rk9u1PHtH/4arL2murxMXC5TmPRxyKZLxMpCtF1CKkicdA51
4F+NUkTEJqDZVeRtjR0pnLFln+VaLV5ob0jmPKAG76TnY6nXz0Pzaq1ynONTMI/BW8LyTnSW+w8B
l48dav3AzBSm0cbOtzoc/naGvKrbZNzd6ImKpHcWXatuNimSHaj6sIWl2fko4WEgTtDsaZQHGvXg
/UhRzUmzVpfvNmlVkI3UePUj3x9bslFQkfPs6C+ZKAHmSLhrGulX+QEMXQFLYBYb5FrTkI+tSa3y
6opwiAPnvBbSFu003KD2h1SO+F24fo7tRlP5yGrobGYwREOUehIbWGOToIzsOqaOAKk/5VRuxNun
CvKB0MoGvwq25otFWvVGByeENGV0Ha7dqwk7TxwD+1kha6to/KtKLt0e0BbLaAWU7k17OX6liDCn
KkTR9DM6l3nR9kLqORUEBoklpcpIIk1MjtUT018abkcAXjoxfQz5IP5IDg7I8EIJk5Dw87G7ic7n
fZqL1xAygDQu9IswILG/XLR3V5ZH297bhOm5T9x+DC2V8mg86vl62aGSjdni4OwdD5EtluvhlpVs
4huuOum4Jcnxg4bSfNnrvV5YD2KzAG/Qrjcshwce7kfbzZfhrjAM5EGD4wrbKeYB9IQ2esoSbcnC
HJYXjeOH2H7sDZ4xPoe0Ij3xinScP4x77QQmImTVi5LCpPnypH1sSXv3z9MGMr6BHiO7iV8ncd+H
ZF/1Mi2rMlD10hx9bcURNxcQtK9YCXBQ/k8pyvbOHkqgme6+ww7BL/DfxUNm09g19n8WatwBac1n
xWrPeOC5lolnrsoU6L5AcRcaSalJpTeIwYXv3oLBHQjqUvSPC+u5l7YIB3Bgt5UjPlov7+homDCm
6KpdfsJIp24YLF1mVMXbLHqP5Zwxqmyx5JzgmPP55yAOy34kCh+QW/iB7YWvz2hlwtan9khexp1P
ATArqI+Wuq1xyQF1gjypVqQQCI2kI23N7My9uscxyReyW4hO1UTulRgswq40rTW9Wo43fNV+GDlg
SuqP4/43aoqCRaUo7V2VszuKhLFcxStxVpa5+ZfP7k+aOOb9FqzQcOEgwe2gGkLwpK0JL6rbj7St
Kd2WLMHMHsc/jJss+nD2suxeyoYIU7pq+/73os87EgCAE5+EKHsIGUxWpBAM2wfuFkNra4shqpN1
n3xDbYJoPSaWdHD0H8flEO1xadYZgGusy6XUAjJs9vES3Bi9Og5zywwiXT8Z5HRHBPDxPNzb6Cht
wimbLQsCAYW+tSfsVwKZ/QSk3qjT3Lmu8i/DWCRGtCderIURDw7fhG+XwtyU/kpzo0j0U9nek4ES
GdRQO54sQ3C6vAsyQp89Z8rDnjR7yQ+8rMyr8jBcjeIAVOnwKnujKbItL/U+2/JRq25jBs+groLS
AYK52PYcIZcK7a7R+i7ZDWNSaVvb/TYUDgTjfBXN3yKraizHHH2HIRC18QCkDr6FpP0Pu7Yzzc0J
B9W3p0oouz/pqWoCGQz07qLaYdTfI0qZ1YTY/+stqlPbLawKUAFmRyYvQbngh+wUjJAxy+2OOu9H
Wk6Dm9T9wkF1smz9M9mVAd9TTkbzYoQniOAxr17GLnV+dDNhepQTzGpOVK7VFTcWnbknK/tW/F5I
qrFF57PHLa+7uAJpN/34Unrs1QTESPrIkkxES0Y8Bdi8tcyh1RSBFcWn3iE22KRrE3YEwTYuny3P
QtSIuzfyY6tNN9AIRdi77PcI+ccVefYLUHE8Nf+cheNhUq7c9zH4Cz/3QF1EKmnYU3iavRRSP4BV
XqhiaBWPMNH6HjCGLA4f2ahEW6nDIjz0itu6D+/4olVkhnTyEshua7fyctoPnG9DekAwtr6aD7bS
Kkcs8Idv5c5Lyhw0n6fqOPIGFoJ3et6vFepRH/xw7k/1hbQ+g/iVqyxl+5ig0gS66yzEZOF13/e4
XB9wFOD6mo/wbA2vVxg6F4zRBREyyXPjsh52hmNy8pDb0EF9Y1ofLHjSAsscJQe1V9BLCcMJ6Xei
bFFv7/hMquH5llwQdV9n+8a3np8J7w/ZcQ8cLBOeN6IOQ5e5HvDkFWHHZTSlYt9/8VtJ8JMsdCmx
rTT3eq5sOVmgxtlcf6ZZGKIzHYBRYHUrZBr4feB/+391FYjMPhZX1HRrvtWMrWrstGV1eWfR1P7R
7R2DxBALxS1SuZEculKfyeyVZ1Rgrxh+5PHD8YxwkcS13WgS8ydUbKq75M/5hdM0bQ/F0em8Q9YA
JMtfIP60DmS1vVjd2XoYzo+HOa0ik07GmYddyqthhHRmZFwi1djUjZsAYhrOgaiOMVh6aH3cjYHQ
BM634BNh8AHzu9EtRlh0B4+7amu9+MYZvp1FOT8RljT27Ll+sBvfh6uK1UEKXvm8/nbc3IRyuAGd
0A/gInxAciS9b+1EG4PRSFYctcFwo2XkNG5N5UNoNgyupwQ8UJtZtOi8AiapVP5ngYpeKVPhM3Ne
vdBNwlnyz0Qlab+o+GGvNnf1q6QmgIUvfaXfnqieJreGxCPcgLh81gXsv9MJ3+YwRDuYX280gEZe
eKYJsUGRDAWXQ19NwkEXO73/NGCcecTXWQPo5bQCX97cY/TZIX7rpPSI2iy87C6KFNNJTmYYvzD5
Oqwvnbd4pMP/ggUabqDeUGjl6dgNc5nXeTXF1gwrQQ5Tpfv+9v7AD4HSDWIBwiymN6jUNj1k1Gkt
HIPqId5xkKI22sFePd4PnCnnPYJRoqrcrPzisBJW7QTwVG7/2l3lOv6rDV0qGRL1g+OTQm7ta/y5
9wZz/PY/k8Uc9nbPzOqW+gr5Hsd1yHUDPCNj8ZH6o4k00zAoZdPklF4TaZEQ+dWUZlfWz5+NEKtE
5akIQ9Lat5uGorTahO3uox4Fen5ltLlZb3K0CV92ElNV+KFbPk5vkYbMcESOXB+7GREVEKMLO2Md
8NUpmf5WriVJbvU/iTcAEY8mUvwJXHqZ93dUX22L+8TM9RqHKPKWMLQCKdbEa093tWeq60EmUfxJ
TFDHbmMt8Y98H83eEIja0s7sqYaMu/B+LDV4z/h4tGsfIUfL8tQRFRBrx/LOeA+cQbyLwTMvg1Hf
XhCUiTESfu94uBPEX2d8Li+z68NRCzWG9WuuSGa2dNkaIwMXatnJnO8LimhVXgqfsxCg5VXHUVfo
PJVF2varCHjuLbM2vPqB53Bb4Ja065iPKgqW+nFNWD1iIWSpJecxLgyGe2VRBjaIdvbp3x0yN1MN
swPGkNrSjgVi1DjfI4YVhO39ePd4tW+qv6e7udPNHQFPM+4iI/rAT5Yz/gOa3LujkDGMPh2OnS2e
DOz4JZ+VohK/lBGyJGMrvQgVh6rzN/+GnHSkF67foaFoUJFdnVFmUJpui9d0BgNKg0HmrQqgGf4g
jr1AYzXtzCa6lltIRUI6BWA+d2JBdauiEEIumY2L2n+jdzqLzhN1tHzfOBgPJavRyQXS8yI2GknU
k6uFyt8DO0Yr4O7CarGKQGuxj0/MfkhUQFPliriyfYiTQMabQK0xNqGZb+tbW+hvArNqg+Loml7T
+L5koz2QoPlZRpEIM2qXy+SVm2XicDqeNT9GY4D2Gyhxrl6cKWME+IZEZTxEjVryUpRjbg9Fj9d3
V2uvtSSngQzIEhE99UlSFzBJGWg4Za2hzNnYVI3m6zxUwe/PiH/s0+nkUdofjmkX1NGHpKjqJkQZ
Lu5NXRfJTAxKPMgjrj2/B50g1xhVpxM5n3HHiaZ/Evka0nRvBfgsd3ivnEIrTfac6BU5DwIlvNr4
AKifk4jkLxo8CgKQ8STJbKF3cjpA/7fl33vcfdwZ5ikXswH2AXS2HPmrkuP+Ry1hCTPccFELkszN
Y8golzVczj1uJxjgF/71TaBzdHHtdgVnfmgaArWSUr0+0UcSKxTEyjMEYTYd26lnFH5/mnqr4bHF
mxcjwjxj21xXJlMc/PszhlTvApCVExU+E2aFlF0gdznQvmm59Gv0FUCQy17tXQl+TZElQKFVS7n4
luF7awD21AcXrt8MlZ4YQLoPWCyqiT1Uzr6EK13RU2IAEOeRdXusWHavGcAL4/usewPXdqcb8w3q
xpzKradQQ9g8054kD4X+gIQb+m+hNc2FsdGUs+GXXArj8c7Wa9ZcsjSk1/CmZpCtAJndbHLZ4ls0
dqfU1fzRM7BxwgfJYzaRRJw0iICRyqEV6psj+rbUDC1g6PlFi9od58fJ3Z5lOB+5pW6WnAl0UhWJ
4S3yiXYIl1g2/yYeoTuXkUwe4AITkKW7Uh+iY9m4xAhXQkWhgQmU+4/nUrQhm6fc2zcpyzBjb3yY
KZc1IO1HhK3gnLkKgwfbKlasmDxrUcd7p+o9bnSbwz26Tnkdg90Xnu022SFH07R3pdieSOFCJdt3
4WhrmnXU47bSGnkRaI6k7Qlnj/I8MBW6WpHEn1qIstZAJyzY2wN//MdkGUf9U0PFknnDrzfOd8gW
lE7Xo//tWEiBxs0KOP8i4ZO4do0Ba2rlMWTG7eKWQaIIe+hR0auMUWIqeRetRxN3bpKVxf7a6yCw
fnCQOjMNMa1fAD2W0+wLN6xJoF/5WdW1252DpMwHb71f0iVf4K1SKCUdoBuK9HMs5fmMI1Elmxnn
ADTkkClNGPfXIlEMfgScXHlzbk1zZP5NBho9k73C4VlMh4REqDFrnx84atimEEH5uEdARFu/k9cZ
RUPLrigRepv2G8NDse1wGkX45qCwMel/Hdn3SKs1imV2o5x+1PiaMgNjZSQ43kTfaPTUOMPJ61qj
M5Vn8DR2LqTXDirUxgUgySUNHNBc85YdsXu3h31Lf87kbjckP2YxRIpepIDCVw777TEnqs6pjEXX
MNPpo4Kz+o1FJmsotTGyDK5l4469O8CzHg8MPZvqtflTlsHuk54ZOWyLIOLC/Oc0FTYLObL6kgw0
e0rTMTQErEYnCYEMJ9hS368KfyDftMJgNt5FP4pHCeyCErqSbx/lAT0xBf2+o2EI9MYpTYlKr7QW
2gef1jiluJ63tihP1I+D1Od5oUjf9q5o/zuyB4FMJV0LVlW+nmM8uDKp9bm2o+ROy6PCpe6cWUxl
d03nCm9GcB9FQBEDUMM4KPLjC9RClv8PpOQXK9dlEw9ChNaDtJ4amF+FaNlhithDn+D5Z9IaxHBM
8BmCsvWJQ/KKnac7WdBlOS74ZC20pFRE7od5NcRA4/zMKTToEyvedXcefHcxk7XsqZB28Ab82wOR
AW2WCJ+F7PqUWeGevNjxDWk4xX9J2QkphXbH13tSZVgvx47yyRBV4uTWHrWxIea61eRlToyaSHFJ
B4RICUacXHMu6hQ8S19Y1S6H5cHxrIFly6SPk2YzC59PdITc/dzzvUPHqGU2f6+rpft18eBHQmVd
brhxoJBsAkk4OL0DXYOTEeXmS2d5xECdFZyn1zfto+dFXd+TlGKnvcDRnAqIpcm1EbPqPnfhOOpv
rLGAPyDbQS0W2dwp0/8zyQpaxc3GhjWgzACt/ve/rQ7CjrzH2DVj9IglL43Z7mTJ4hafROGrVMYx
ichuH4CHR/yK1Xi3E5TdOROCBjwOfvNh3BdMAw8A0kIEMihHHlqfZo7l0lBLTriKprBwKikyzi4T
yrLtwL/WE2add9C6eCqCZTgOuPvi29kDby62wyDVZXUaHD/98L8zMgZL9yNG0VyGeI9PpaatfTM/
YG7VyamDVviN751JPZO/+8TqVRTXV03BiLqmETRSChCX2iqHjj61HarpyBThNgAEn1GNhz0wAcKr
HQTqgpTpnTa+9w99wkUDO679b0TBo8pzzqDt3HmgYcTUS7nA1XnzQ40FJrw5BgfWK31BIuhtkKCx
wati0tLbPcjqFs/IrZ3LNpH91TkbvhgrtTr6n8J/oiSRWVm10Z+HzCpBHXT9TG/Xfa4tU2iXj6Mz
0q5lAXvaJtBMwKfJoGuh/slnz2XRA2GizXWZpHkmNij2GiGHX+9es5LyEtqmHCQJbdS7LsRBE/71
fYqw5+GzotnkdnUBGwzf8ZbSUD5gbU+UWg0SywACJvLs7HP/sNF+FkdnkePadZAViucDYITzWdBw
M20HWpBecqWaI9X7A9iTTYErOnY/+wAcEAmZ+YXIgmwjys+pYr3BrbbOQmVJwkXcv0AddsEUO/2k
lXBLPHPyVHwsaH06iAqCge+EfnRFL4Vmw8JE9AMAdE6g9ZIPnQXdLcjGLwEZRbeHJnDvh3Nlqj5G
tHxkB9QfRjvFDFXhah8mKFZDGfuEd5EU9f2h6am3nnw01rRWA77Ly9WC/jY0/Xxrfnrr1t2bBofA
NdkVzwAIBhoxth2Yyoz8PngVdmjENp+8McUSDdPkybX2fxfIELgeU2rObafO1SolXh17GzlA99zq
GiJw96DPUW94zA8g+ZbXyo++ur+PEdKRac9yZxysHcy+rFOjri5ppvW7/jsxuC7lqWGFDb+itcfk
8zQpGkGWUf45mvbpqCEYK8X8GmfeGW7sEIj3cobIOIyiRM28nJNap9iMRSjcnG099zJmuBFCdRHv
N0GFGK4p29d8RxIdD4pfbDJ9qte6u3YaGygP86tnHB5+yVI1kKSsuxjr2bci1tgtN4csliggvmjv
WiBKvTyBrUSYJZZY8lEXjRzxRSYrfJQPv1BWAbXSpio+unboCX8s+1EoQ2T7ZuJPUgQjIqLQrUxP
I4tPDe3l2MbqJCzJi/6YOTQnqKt944cEM1TjdPLdpAC0fRsROqdNQSvE/csoefnhmOVsEfKQnMuJ
+9wvBA8TA708yutvfMw/l8H5/elh4PKj30yoVTFTIvi4bFMACN5jNj9fZBeUmIp9RrICzIB5bTcp
GDNJDeWQWEzPh0is3fqlpV4nKOveDycQZ88RaTsVkwhDBNTD7ptdKJHjB2zoKSR+N/UHRWO4DkTd
3oCGZlLBshgKIxchXk3mlfJdiqtC2HswhU9pniznzRb8RsopTw9OyiSu9K9of2z2s3fIspP/GN5M
08IjPSadOKEkYCxH3+C1svsOIoqlK+zuajC2Db6gSdiaSIVJT8B1q02K//n00JI9bak/IR/jZN9Q
BkkKscxt2rqyk/RM9jwCqgONRsg6PPoK+Ng31uhqhdmdIrAVzITBDhH42YlnPWnhyKsYjmgQQ11d
noDjdc/XkWJ9893Pqb2reS5Q+zRqvX3jfWn87FXY8vgE3W1z3avvIL8eVW8qKcRsGWTQ95g2PmGi
Fs3RniIf3insZz1ImaYYqidzJCtksnPMug59RfHb4GkY5be6ED1Nf/CIfMlII43KEW+jkWQLBKGq
KnWeuHLAmEiQ4EiZmrjEa3q+lKCHAs4HoXKeRheQEHavHmPiAEiQED/bqs5Ht4+H7DjlHQshEOWc
g5Q2+jhIaM+p7PP3JrQtT19oswcBlm5uZHKWq4dyfT4D2kOybNfLi9XM5lXXBx1Gkjff2t/FSczD
wZmhFHTq47yhhcASSbGeY0xGmxqDZ2KVlmwE/eqgTngc9pAkNpwAUvp642UhCRULdP2Fmp7b+UGO
RpQu5bi35IcFxS4pWUeWqqlRBKCaW8IAPfvXrQhD/OGGop/pXJraxCmNr5IycvabKCFFnVYp8TBz
1gjE25GojNwjKXwkZJTLGpLhmhqq96lhaOdsecQD/YR1J107zcgrW7bKsERmYErP48klx08OwW8s
u679QkKiqPC8b4hmfI9cDbsoGfl6HBmaCLejGlBDHm0wPkfv1G3R03/d+MpWvXZqiG5fQEDGct8E
X9/8kdTYLiNbJ0z1k7MBoh6SyKJzwOZ9j1TzSHwidbfnpLk7jVh+GpAYsnxFQTiFSYmtMhsOXaiY
djO+E4TDyAYwdnIKff0+C66V8n/UMpfzdHg/8C5/nzSXvmEzK3YFpMUtrUrkk52PHxNNEcGKH9ws
aLNsviJg4qM4vkYY9kNHzl4WcsLy2Ns9dWS5CFqwMpEt9p+T+oA6Q9KIF0R603APKHq8TzkgMVQW
qa5w7/uhPq1fUnD/OCJjFJL+aO9kEaCwJOyHrkhnuJIAn9TRKTPBAE4I3Mtu2huAh46l4SoJEwCq
oDYXneKARy7JKFpNiVfN3DqT6IPQs0xIj/4ojscahckONZ7D+ULzCC3PR7s8EswKn5VuDRmDwGkn
neixaL4fng+KOpfC2ezRu4BCxwFcwjmsT2iYgWo/1r18WauQgiNP2esB2/tHpnBKin9p8ICdmhyB
dWnHBOqqlsly8/MwDG0AOVGYonhMvmlFiervZQNzLoCI/JQOCgCxV+SItVdRqZvqRLeM8HdEAec3
g1+WQJVIO7ByoQgQnESCMAuFoUKA5t/fP6xb5BwY+wRbV3BNUD0Sv9qqDx9ntMReL1lAiLtXbsC7
aIelYHH3pmfVa1ISbGpDEVaz3mip0G4XVBfHMPuRLEBJIbQhwSi4clwngjF64JpzZjRVb03al7fA
36ZRCIxSs5LAX2b9n2O2WItBqZMZ7eQt/zbLE+GivkNP4ejP/SvRpHesH/8Mozf9PqMyIekPCYAP
nlbNF4weUJl7wNQamEoHPbWIxn+6n8gQ2tKwoSaNHEoJn2pMwp5MDgdY0dmVM9xy5By3klhR8Jfp
YH254oKshpO++GAKfFHZr3PmaC2/yfFQSv+gijBdpXfWcyYKeYJC4HHqFIsqmg4fJCu7HZ8qSFEl
YP86eD3ifhkUNvnipqHsE0lL8SYmEs50BGQy6Hzt6GxlolKu/dblAS/76aCM5kAL0mC80+pFpe2B
u3N23EcFYQtYvpQ+Qd6v8Yzs5U9Nn2cCowlw+6or/HzuIlTffaG4Bia7fb6tpuxDu/TkKSBNExvg
sNbx5c1Tor09hoNmAzKVgHC/8Oh44vDvjoljj7HpdnxoR1lOD9mofMI+Y/+F2hL5igluvleRv8A2
zpmjAz6esMVrsyuVdVuZItR7Cmn8UbhszuloUiBbQr6xSGkh9VL31svf85fYcq8kxfuDJDvGsBFC
xX3+gc/WTvLiuQrBW5eGB0K0Sv6GJG/ZzRVqLnJnGUC2WiAEkR3MYYLk1OsGhr3iHULgIrVr205t
aTj2I7ByXzMcQ7ypypB6zpBa/o9AgiIKoNhWdACD60tL2DA8pJgn6JKqVDub1hg0EUqfluj2hH4w
zysxb/jCxyhvCl4is2nzUtmKn45PgtjBvO9Sl9AoX8+teN0neGJh1sUJCEA89btS6mRJuIHP9TAk
jZzjyC02H1j0XS4TSsd5Fpl1SPtV1irc23I37sd0vs7hO+JR3cMVpRYCaUTYIDbK46OhvjaXJ26v
ixTbvOWxSBeTO4H2obly9sF2Wcviwcm0z7U7/va41MP/kPh2mI5NAAcxFYwT2YlDf1kFrhAM5po1
AVgufn1JH92bJmi8nidCHcBqvsFoile6EnPu079THqdTQX3Xj8SPpR0ZYDAOIdkmY3zjFUctWOG7
dEbnq74FfAgGZ41KwfOtASolySVeqKKCJFpCqmaqHEZ8svyg5yT9lpFzSnK9ZABRhMlOiNQuXxS1
pEQmbPZecxUo60L0XdNf5VL9ZjqEh0HEkUEERKWt0lQdj+3FBA0A2gIc92Yf29pImudkBd/P/DCX
PfDM3YetNjjBc25Iru2sBJ0AXtx/H7ttAMmOiRoitulz3aKSwv3DHRFmkQZbtEzL/juVZJLarrMt
5eXahd2TLzptFiOjESPcxyNYD28v/TdJ0EI2Ts+SZ4SaYUjofQ+Ar+h/pcRO7RFkIzMoQHxpIWVa
9o8oUnfnfZjQwdpTBUxMCB+3JlQN4GnwHahhdgQOYd0Is1fmNCranjgSQbqR70hxXmfeqtpz81wa
riXJojWqnUIbICk2WmkAUCGTOX4XKAJFBuVWyOHdYwxSIUrhxBar64J16wu4dKDcbBlfIqShs62S
lF2/NFQCrYFjNX59kWhB4+SmGG337Om+EICzDIxCb9Jk+AcEVoUX68VHAh8yi5hhbg+177oF2sA7
4xrI2UC22hCA6ZxC0OBUqGs3Rh5Nv7HiWLEZdBwNmrDy+viJVtfDntwaRDQYpr5o9N9vywvzH7bz
xRXDsgtzLpP9HVkvHlnZcVb4t8TU8mengWLgOqfWvrNCiRrk++ZDIrUmHZsZFFy5pOfG7NEVDBfX
Z60OsPCMcBeyXnFbvav9g6R3rsa5O2BriX0SlXVLzA+jOw5lRpZyv9rDWIBJOcjUrOEouk6ucEJr
iWm5UDEAdBUZm2lx/OWTxghfCbDV/sjIygOMP6uMrSPXp5GVUNYffhSyskqJi3czj+2vl3/rl4YX
lvea5qQrXTA2fDOEeJpn4gtGqofBPV4CvD63vIIO5XWlQ0RDYLCuJ91pR940nsz0imoliYhqG905
C8IDHXvu6vrqLvWiyTggaMJywVZtEsTzFjaHfaSqBBeuttdMp6gBcSgwvmJIfF4z1jSZKzf5FbCd
PY+/MaRseKFtOdJ6/lKHacy0C4LRwkx5uE/Fk8K39Xc2Uc7bXauPtGi7nZSP5jFPdZrLBsNLFCkh
EhUXAi1R0OmSt0Lre5YZgUr7+smo1iVkA4nv/DzmvaGwqhj6mWRK52vuxdOWnEdc8dJj/MEbSJjs
gRgpPxI/GERspMhpq4xH7kJVGOZNnMb4B4Sn/M6IedVOrKEgs4khEm8mkOdyJMxCeRIJCOSf3BSN
XnWQlVfbN0It3vtUyUIuif7ASWDsaiXDNg2svwzLA1Fgm187KfPiWMJCMtMYTK/iOm+tNhm94Y2U
jcWjkCAcWBhaf6by30J2lIXUAOi181CZolzWA/ovA6jRaw80CJ4gmGnzG9eGzBHCDeKWGia/04VS
iD1TOFgjDlyxlrGKC0aDHc577rfgMskk4yH0siU53lyBZ5wJAhoCZmkzZu/bLxr7haGYrASepU+z
MrX3ePofOQT8YB+BvW7Jc1ty8yVnJa82YthsCZ+gueDdATdHgkWGcR0rrmjaYdZQOAZpOfhjP+py
eCmEe6NjYpvxqFp3OtQTK20P6D3jhkjdBKJtL0SYLqztBLOovjsGHHzccZTTb+/1bNyu+HHOsI6m
5Thxue2Hw70dktNDJwSVy9lR+rJdf55sh1E/mAaui+JBkvg9pnqHYiFMKDzNURc8jKLdBBMH/IhB
UzzZXdEu5TmRDETBYz4Il4lwHlm4Am70DehVT7NPPkdCXCoJ3Sb1SXhcvrMbZrNoCB1naFbWifpU
6WT+NOecsXDzny6gfQy6YKdnslZxVjFRgzp6ZZlKzZ4n8poRNQSLVIWb77XVs++zHGhu7mRqjHTD
/6cK4mKC0S7xGqPRQZqg2wDZfk7IvnWNhTTLkNoe7DEuf//n5mBZIpv9+8iZZU9W3yalcmUG57PF
d2pWzXlZuugU7UMHKF+2icOsay80lUxKlNWci0+WqNBlG+ZqOkAQRSb8S9Kt0x1EP8a/9pHSgwXM
X0FqfMI3Tu8tD6H/fsYHfb9ekvI9NYeQvdyWGwzdGqbGVuMY1etCu5IRTwssSz92EtiNo4RzEq0z
ZDIaFKG1j4P9G+GD+9wvHbXpw+f+nXT3Uey3PgVNYMDPAUcM7siQOohZBaQYRoAwQ6RGDogqen+P
C0Kc0DXTw/SWsk98bzdkfo54f9h3pybL6m8BKVUAMLoGt291zLPBQvC3/56MesYu8rCfEtgcWXhN
F4SIF2g9ae2lWYvAMT/owFKylgROZRsJM5rt90H8r5GNcTfz5zB8z4NB2DxlkxaZDUIZTfz/G4mZ
aw81vOJB8u1dnZAfazVl975NpqY/5L7uxXAHAiW4ZAWnGo3Ob+4Ic+ytp/3GLA22v6OP42FtlP84
O0QLhSJtGnFIK6DP8HgrsMd8KW7NIyG4iZVURvaQvwb0ndTkj0oO5yjUrQk+fR96aTfpZbYtzrff
4ExRqyb9R6oc+IXSq/wIe81lm+ki/NnawlV4e+JORoCxu8NELNCdizPHBKcyElOV6C3w/nwcTneJ
P96IIeNYzPCbUrKzNH8/8XymXSPxKp6TBEq5kbgFpnvC8cn0Oi1pUtekAWzDbbGAvV4qlQNSdqws
CUbanB1d84ICQbNV5woWLQqXg6KGUH5vFMHy4A3tIGYy9ZAj/j3daVTLc5J0StDHxT/HNaA4CcQu
rzPrI8dwZXhwQMXMtJOwuuLZw2ulV5dw/4b3Jb1PJv6QZkTFp9+gW9i62pY2isSiXtC2m0uIwplk
QhS8Z3QyUnEAjJMoxinIPuTitT1wLvbNwktQ3JgXiKESniF42s3oJ+bfjq5KHaPbxLrQKJ5V1Q+3
o0Damwmg+NhcswGIu0yqK1Ehq9gaZX7Bnt+0Kb3P0nownFXvMhFlj76hbbBc2Mw/bkOuhE8xmysq
HYhkzMQYMnoJV1EYSd1zp+ejGrHpHtMQaC2rpUwys+VQkB8T5NIFHd+KCWD4sTEFVswnbzm7lHli
NqwP9qqd0mLfN7UJv8d49P86JStg13I3jvhhsoryF3qEpPBx0bEZ83ckD8jaEXDTh/MhwIsi5Pex
2J1aNOo10UUEt4p19+xCVZ8Uu8lnh9WoNC0ozp4qpy5znr5vAaRD/wEhkQJ7dYPbFwCLxAkLWbRp
a2w3PR4h46eEcjl9mjjydihUveTfGO9S56ueNI1/B1P/K1VDopCdG0QdD3M15XuscbTf/ytCFGHC
NSXwYlcA5yl2D+24Y1xVQEvVJuUtBdN4uZdHGkFtlEQ1MKvchIyUm/+t06/jdvBgs6QZ6QoL0PXT
yRlOUMcczESRaqXXIYN+dgM/xpfgSWYWXHVKbyrhOHSPZkhfDNWJukliJikPEPdM1LHI6KtKMy1R
MGNXrRbYi0OGa+xJBJjMUlsamno4hs4VXbkwpN3l51kbiuHH5zhngY4mF/1PpnmkYNMyNnf0fYsY
Fo7IGTbV5yufimw9276fGxsdQAez+DxRoCcb4Lxi4K6LTDwB52KTaltxxbl+Y5Hi41l7lMUk4A5F
bjDpJU+pGIQasDUCzG5aC3tkp+vmwbtxkwbaxeqEyBABOGv8LN7p0kk+zOXjMYprTz360seuscp+
XOmP+1y/2Q6cjC2czbBR7N6F+napAFZWvbtWj02RGUhnVrpRBrhctWXv5cgjvxY+DhV+ZuJNFGtN
4ph1Pok6w2/PPqDTWunHUEAkhPbc5tOvNosmD8qQjZ5ygmr1aTiqLiex2TDWalPrBXi8jCpq3wHv
TAoSMzjWfZBBARPxVKDZcYP/7yXxwz+61yiw2pNV/vDhXA/gK6R7nP6cdZD6AMNtwEzR/HTguphE
tsWxovxzHKdzssfpbsyaJxA5BSG6PoA0GnJTJQg1V5kBKbyQM3CLm/uQAi1hOf1HLPSBwPmLDPQZ
gThiQWose+tCr2V8FuezXZj78/gbaHXbgLoMHMA4yLIDwA/qXqR2a31RKzYhh+puKAdF1G6RcNUm
+0y8h+pgNVGurrmKZZzREbH6GWrHA5HRlhQyP8Ab3BwqNEgaiPVix3fQaJWhL6h7q2OIUVY2tJ34
eLMHP/uBr2GFc2dRBiLZbGpayJ4oxkdUoting9X7dVtl69bubtUobjjoeiUmy3H4iIvUsnWEwZFv
GS/8/p3XILe1ddhk9qRuIZv3ZC2R39jKWtakQsROOR18D9+bdSzhFzJ2I/NWAkM9830Htjp3IqZ6
9QaHI7NSpNm2aG+6KBRV9GEQ0bVlsUvDjIzBE9R3fsypcUwqcywPLW9W9HMdzEoA9axkjcIdBQrX
rSWLvu7hm71XmkZLBKlwTbNTwWiNIfilYdZRm9soXW7Ve07gW35cbTol8AP1AHEPiUXia7tigAJ+
UWQtY24yV7lGo3mE9GLKl8+Tp9H1LT+tz/tBooZyJY9XXk3zj1ke97wgE9Yl9VaTYoKLC85ldvae
HKUOwkJfAAxiLTvm/CXiNfworvyeHySgTdegJENghEJus+NcqOE886NgppU7Ifx/3ekqBgOCuQko
wFXw+t0nluhv1f5cyk+Ezitg2o3yhp0QWIV9huqTJxEHZyrl1e47Tesh96aqO3gBJohZyzXlvj2x
ubvz9ZzDzkaoYbik8Shcecm3fJz9ClCVwFF8CHV4l2V2m6bDhx6ZBh2smgvGugBgM/hAidt1/Et6
x+lE+D5KV0NWyrE5wIF8zi75HOcCyUWUbeZEJ9cMo4eflzi2KgaJS0ektsxY4FR/DCJPFIISPIDR
S6EvGAKoaK7FeVZFoMfyyfy5Iqr79QkkkS5nO6Estg9hEOFTtuuqQO12OoSdu0lx4NfzqJCmFXhW
eJj8HmL8pw9CmVToZfXWimZLLlCzkusAoE6FkTGBx+oU2E1qFF3NMvkxz5ivkHnrvF9mkLnH3r/i
U7+5SVN1Ok0FliGbJE4Ux0y8Seg9LvGRuaNBr7Bl2oWNqLCo4gC0bsuVmFlo+3q54ps1J0ldKjAG
ZUB5XyvDZnNsZDB8RYi2M+MeP4yJ7T73A3BQOvmyx+8g1VgEzoVTOwbScD5aIrxR8i3w7+17vUZ8
b5KWVY6UrThz7aZWpBl4irHV8TrAJq11/zt4guGYTUm86uJTg+bov1NFYKTr1qrnCim+Rh/Ynuy4
BQ3wlhSvdCV1h2+GvMd/33ISW16NFNmFgI8pW+r7RwTjxkMJ37q/+RKDIO8dry+/kM/Zyk3wBNqf
xZDEH6Vu/285f8hs8g2slA6Zp7BpVv/cEWT32uEolSiifF1uSmi4Lka5FRIp7xnO8tzfoh8Ktg4E
/TakxopuWbdNTVUew37e8jQTfRb+y3EQ5m7dJQyYtQspiQne6EDQJc1hf852CPqyT8YerM57Zlaf
+l/AOOI+4AWLzfXhQEcwqowgnN9oiPoduXeifLkW7gzUfKfzv2p4/umEFc6Fti/tRBLzYjAdjIqs
stcQjvOOLR8/Z45zlj6R4YYNgH5tm8upEioQC+dlNC2pzYQxhUv8FOeQU3hh+2KsdyKOuzoc3OHo
miDMQvKbSC2J1XUOoeLRwoRHRFtiJeI+h4B23Xk801sdmpKYPUI5Lp9v14eEwPkOMH8N3DGedIM9
IZPrbKmJf0MapWQox0BoIA1GGJz1b9VNZ3xehCf+6GmZHXp43Wz5yRq38ilim4JcyXnoSM2f8QHH
bXqbECBH4U6hrp0ousWm/2ViXstOekMwpwjvP2GYmOmtVY1ZLbtaLuI/OGCfXo80inHPofBHL8eM
lzImlwii00/IX4lfDDCC6NpK6RMOlKxf/qaauD1mFyHKg9pAmYVYxzswBJx6C9aunV8Bvv/wOJWq
mHWxLbDPoGSRKqZrfRlqAyB5FZmKCDrw0OMDF2kHnND10GYcWE6alSbm6uH/Tz+TMLNyJb+4ohOQ
3KI38Xlm+Sg2Bs8bnoX0E+ydDhowcHSjptOSVHhccKMb96kShSfDw5skFMosEEgUNONLmLoHxdCm
dpOqUUHYeSl07Y/ULnf3unu5oEGv85pF4V5kvcIGqqMuqzsRE7Yi7lk44spvQ36I2gASuc6DsV7d
5n8Xo0W7Zm4tsVN3x48+/k11u7W5uZqaZd8fWxVjZfJSs+jAoSdUR4TCsLtHNoyrfss/TcwQbkyp
NAnLXLnlXFoEFnmMLLrX1Y3hm9vipZ9b1O+MMKHpQbQRHLdxxU/T6L4hoOhrwtITw1NTk4W2thHW
CETq/xkqNwaRPXFDz/ZyHLENPSjVkqFbBimwN+16BHSPtL8BN7aC97NnLQXDLd/TGVMNkdI5jYNa
vs5ZZNqwMG3DUiCI5tCF5k/igLvigkdsRhazv1dR6NIvDIkasf+EHRa6BErcpgB9s94QuNZ4zdMr
bA/5eE6XsjtCbhEayEH1Q8nVrJsHHqC909a5QnqHtL6s4uK3qnWMPSEYhTv/AxgkNUGAcyFmmEZo
MEtVO4xlInjLj2psPVuxVWl+sUjTldxYG28zuNWenTtZjsr0VoSdaKBFqeg6dPFjIaxIMXYGauPw
0U1NUz9Uq2fzAB/cItnHwCJvvSQxuymduHeGh/IlRlbzwIklPibYURYXCG6Kv58bFGS/imPTxA41
xPwp7OzOk/4lS6OJ0JaBA+FJH4DPFKXz/Zig3CF4d1tvNulfsHL1KnpYgsg7mLZ3vhEd/vgwvEU3
6ZjqtBrRstEpN853fZZuMHM6jJqIAiW7zfSkGFYsJyU8B3Bt5Vp0glADX6CMxJlXyCZgc49OcGvb
7dY/XN8DFIjFq6Mj7Z4GLpT45nMyRvJDdA18/JyTJpZsLZqObjR6jGMH7L6ZXPFlnD0f/vK1K+T0
X7aI2e043yueR1SGfvdEVhhZ0MGdPgqNOXVOT2o8cczdMWE35ZuwQBNX8cqWSl3j5zgmV9Fg1D5X
Ajpz+DB5YIC64WH7B+NKkY3tygG+IPT/YD0TffgkO+dopg67qoXr7ZCzZwrR0moDUm9P2cVwRtYr
h6G0LY8pOQJIDzdzGUCyAJPxji3CTHe7yfK/sKYTa3iPwNhVypSh/SGhE8YfvbdUyy7qy/qvOgzP
/xZEdmi2G948VnO+Ca1UdSEHBS7N5lOkxO1UfkFRihlwlTaU2Zw6X3acfMGrAiqbCJ+Hki0OO9/T
9o4T9yI16WoBJbOiEHyWbj9x+LcoPujkvM5Ih0YxVCRwaBhdV3kYVk3JgDArSIigKs0JTi7WAHNv
OE84YyYGF0r2u7qm1S457CIl5TEVv0xY/es2l4T8K4cve/rTqsFJTDxwxlvz3beUUxEif03Moi8K
C/iH4xhvqYiX2ut950In3pKFZbmddDZAKSvuoArlhauCdeDoc3+OiwTS00o91Vh0hZ0wxGFDJkHM
lxk5vAoEODmDfzLnNxlLdQWq5YdB4qy6/hx052Sn47McV3iaDLXNnntcTxHtf8xt/03tnsC3G7A/
oLqA/oJwFM6iGkv5rw4HE4UYNozDV5yodkzC09dmk478FrzkIIlRwVp0I5fW68gcRUfmxg7IW8yB
QyCeoVTh0jtEdfSlp8h0hoYBYwTrSj3OPhERXJL7fkEYQlXzjUDQFqMME/XEfsOG29W+by9gyOe4
jmPi73mZ92iqmvmwwA0nFULfEjgTW2iFDMasmcg/qOhDJyzyAvaEWSWPLrxK9Kq9nbUcgMHeFvQ+
fc+AD8YMx/tbZcWBa8j1xpFyJAGm37HG8ixjpKPkKy8dtOjb1B40YYvivXhpCC5c5r/i+j91XDFI
yHceRQtL4QACD9C3ypHFq03UzOYqtuZvh/B4wImfF6Yo5keZpIX2yF0JfsusxeHDiSoNu24KXAgB
FZLfcarX0Bkrn7NlMChHvFHN54wgu97hhQFE4Hi/mjLy9CBc9Xq0GfDhnrkpjQ9+DzdHi1nctuuz
1JEATObm6JF+Ucr1+OtkFsofNjGkxsv5oV8APR5CtqkMLuuZ8UeTkYJ12nmWOVVp6ExYzz+Ne4LW
TIo2qqo8hk/uaDYo1j8vcevNnBprdAneHi7tR/ZPS72CPuD0/fHbq49xlBLd8AOcdzUnxXAb3vdR
o4huf4/347KV9p6Ypsi7o94bgTiVD9tOrbiUTy+5I+6KHdHXu2kNq2gUcHmm3R26YsTAH1Q02Wct
gfXFosuKioFlA93WH+zq1DxPrLB8WvgsfJABQzc17cJnd2V5O2Wgto2lra37Vr//lY+LdNHprQVZ
dODxQ0fkap/Rx8Htn2t81uIuyN/nsz1PFTcIU+KyrBFQ3G4A34MyJuQedKrsj67l73LXe4ReV3wZ
r5QUXaaUb9U4xa4xa+HPhB980g01QZimNLHwiNe5DrrfZQV97RdzSl3Ht40SKonmrhVeoXPC+sXR
C9gPsKyOEvAFrAAVSYi2M5FUcMwAP4bVbtx78ku+U4Kf74FP3B8dCsBddKO/9VMXKH3AjAJRc+C6
sjoLSGy/JTdi1G05WmWBQxZ4tToZuPOPZA8qmWwSjFIVA5zJUzT+36JQQmkkh7HPGnkYj3iggL0r
g1Z0Yr+HlcOb7Coa0rqd6A99HNqbJmna/ODeNLOPBHv1KKPyQIdE5buzausBDQhDHgfTAsKSVUBl
Djtr7Q05rU4DeDmJd3ccYC4BUBusJAoaKIJW+Z62RcqfeC+zI8LWIHUpawXF1uxwZ8enWnOFxnNa
1bdpPyb/dI34BEQ5zWrnDBgR0kYYoQB1NjJ/WIuW/nLYo5vy2Q3zikj9OfTe98mPLXLvP0/KCiAs
KQeUnHxOKFEMxFgo8KeRqhT699R625iEUNBsGCcSGLbxsFaCtCf53t46vteKKgJAc/EgOeEuXoEe
O6io3mX9uHb04tfXX7zw0gtQ3O6ivVNZ+MJvesgVlkuegLHnehFv7NMYG3Qira0LFzJ3TQ6Q/WzY
AoGsRRBqZIwljrYwOF8WbiNhcwA4G0GYQj8G4HCE6q/x8mA45VPwoz4EG+g2gjugj8ZrnLt3cpe+
3EJjlaNVtHC8Jky6W5mzIfwjpRMUcYaqmhd0ujWqQECvmqXThf4KFm8uhcfCXHx7M+p8XhGrReVk
LV5dwEZXJmGo6uO7aXrz0hREErWIz0r/VB5xEihf6rDrXAsc9KpiK2g5g08+UH70KzbOqGTHCBWf
jTSdK0tSPQ4Q19YHbATZuC4eEthLyMDBA6eYbFxTEAhnOdUyAK9izJpytzMVTeCtyDbA1GrTynbi
7anV+qsx2/CYYRtJ2uutrlh2NX86qsqTMzOETF2KedMtjE5ZV46pR5WoczxF8C25pVVKbDkQ86Dm
vn9mDBKUIbQmBXHVUoTKEL1+sRuojHLofCGZOGEcHPQYxvgvuw42p4WYwcGMGP2yuqX088aseD0b
jorlo4iTZPKIF0b0MGhYItKRSd3QeU+wgTFljljcq5JWeZPVotWFsN259JvmwH7NNsn5RxaJoJ5s
RHqV8u8tmOou3jNCYzWmk+0wSm5h+CDtavYhvtz6g/8CR7sqSLFaLBdy5gWH6TOnZXkS9Eu2bMCu
6nr07MU2LuTw0eXXuBNsUiQybXFO9N8UBgXjCnxTcT3omBejmKxE020QTpA56kDvZDwL8+XScVRL
Dev1XroHC8MQQMx/pUW/1zOImOgjukLyQU+xVGFsMYbc6o2uH4eodpJktdUIIn0dAdyiLp8g4Vt2
gbbUlT13SN/kA+omRdSPUMJqaf7Q+lgYtyYJ+vY1w1AKoRawawLZ7PDTzphfX6b+Jse2A5UYvHdx
ngadtgokNJFza5XVa2DEN4kP+aZN9OpMMr2I8i9B8vZB7ornUphnOVSicTAIIIdMEYtMgzCdDWnY
yB8vh4RZmhUP3Va3yMesrT/b6uXRDjmqNhAfo2yivufe0Kj0uCco0f4+KQ2FxgP9Tg2Ov3gOtyXz
uPuEehVayLNnXcdtrhsP9qXkq9730VCD4jjWdRGSDr4elhlrNig9i4/ni/P/r0jVb4hJFKrl9NeA
p/7xPVDa3K4wd/ULoKZEgrkfdWzkNBVRKT+t1ol+epgAmqh40mVaFEZyXW/92u14NVw9xQOG+haf
4NEfapBBFh5sP8RIHYWy074nohbPGwjUS11Gc5ywQWcqBadpLikJ4LMqRCy+IamH6+UVqMwWvhlI
HZSJkHNTh53/bHMB+PzHOmb9ixoxkxAK14/vn7tOMtIy8yDPVf1CvYvmdOv+vkgtObunQFGmNH7d
BW0YAATNVoc1z2LfyMMxZ3XS1LIaXW97xxEhA+3EtDtIaAJ/RnzEBmt58JusFsy+MsNxK+fu2qFx
5mD932AuEL2Pv9wKy+H86jV1AnIiB8Jhw6KUZhRVlnD+C3XI1uVova4bo4jO6CIO54BwwlnZtFHa
K8rI7UxF6y77eBok5mqt8qy4KOYvVxs1AvKkqL0OzyVsBR4G69yVdiblikTirXOj/Y3UhyswNmSa
pofAeVKW97PIjNSpoSG/kP9VnvcFLQAwAtkbBY1H3vmaTr40RneUxQA5EssSv9pAfYCXb13SDsJD
DA66/TN06rpA6WcpQW40N3jnwm9JxZNm0oUYySh/RAn5RfhJFhfxO/TaRgpF0gheZ+nJaj2bQpyn
zncR9fyqe4K1sOtv84D5V/6YcBbfJM/nvxXO9uJlHFSh9rQMUg8IgnU8vh2rcPgzbf07PIff1PFE
EB3waRua/Gn6EywfPxVsf+PDrTauGDyN8vHsl+TFGhprKWA2XnIaPuacZxqPqHOlLPZmuA8SByC4
T914qOKB9AVrDhvDqLKoVhmt5WOfQDcKX62VXQ6lG2l0vT8fJb3SCOmrFpxomk2UiXoutYcYyGn8
t1xOr4rUzJJtXSqIWy0EO4ucm6a7TadnFhvGukm/peUPvh+IWy+zX1NRuZi1f3XCY2BT0NTDR9yi
aLoChmaSbx4ApQdAST3E7bJdOn3qSbG+q7Ey9oZY230S0Gaik7BcUXy0b+EnJsafgCx1myl/ZuIs
fgdTlL56MF/0U+qAIMuBvHJurdVLBqzWbgVK3H9xEtyw4GIqmyq2vPZ/NVjICyiezqLeOtLf5V+5
z7ePSoMPa3ARRt0ywozfxRyzV41S9ZAwRBPuDbVzrjHdBCAuXLGsCpFAPuUxDZV/r+3gy4DJqPK3
rjFtE0b7Q+LnRp85xwRzcRqCqh1pJeRWZ5wdu0p7k/v828PzA3/lIOrE7ARCZYfa0y0KUsEK9j9l
62vzDPySgFHRo4TwZnQxZZE8SJPDk7e9OUiAPn32OvENUn9JWkkvMfzK1wVNXgf9WznCl1+L5Mv4
sDcS06sO+9eMuLcVQ+rrI0geZGqSMZwTQnX4g5D0vagys14p12fEhhdBCdD+vlH0jW4+99b5hDpN
5hdVgvZfLP6yZFPnK2sFgPqBjf1QAar3SYRXH8bWqPeK4R9Kr4XmZ0TaoFs28HWTMQS+XgoQuzn/
eu3aVGA8JGOZM0xs4LWRVjDfYsIHMm4ruuaa+9Lr+/eIaFiRDqM3aW536RP1H0cEi8xY++05OiZJ
NtMTf+NrYicLQ3+XHJxStt/jiESCa8saLE8AsPSpz0KhosgPk2rI4ysNaN5kBI71SyQhooekDydS
aFN3CuJtndqAnjrrR/qzSL/4wtUhCbUuhYoOsvGa9tHZoJhep3f0C6Z+Jamdujx5JDei2QnD0b7h
ztnhXP74qE4hRDmxvWwt/u+hoc24BWvQZp6DOhQzJUbE4ElhcU4su0vXxSNFzUI2mpd/8CExKNgm
HRdVHEXbkRpMLZn/ADAJMoTMhvRMdhBZgkROce29HzWRCj/oqxO19gGsVyLRDkmMBGxxj3gUXUw5
AQEfm+8kmtUW/5UU7//eVR2sixtsaqp2XA3T0gw1gE3xbT4+cEWyN8PTNQKVHJRbY7xo1fmEsg3I
FSeqFPl3heGsLz9wKeEMvJx59VhKDaHK1GRnkIV45fCzyULKyHSblls3VK/rJhHeTSv0lDyVX2aC
fA5YNJp0sbaiWX8FIJdaDUc0/tlCtKkY1ueU/MFKDswiG8+v7jk9RUodrHZ1jVGl7VTRAQVlv6d5
Tr1zL3pFppzGeoOzesPs+JddUerCP45uEKnMA96Gezr2PuSivPfE8hGleEwyD8GoKIFzkOc6bvy3
P8e+Gbaz5w813vG7YCgIuWqXhYQ5GeW7v5OiHX4JTcPekIHqFvAHdyEF9c7RpcNj8CJ25YXepPjK
++zRSMAqUavomuF+QfpAVOjtp4uMmHeKxfVZeZ7YiYl5JPUPyX4Es1ISQ0iLhYUXkkFyfgDQIiir
BNU04N6IDt3v5qUUi/uaFyQ7GZEuGq6HD6kil3os3793hBaddDMj0boFEo1Y5QMSU2QEZLwV7fDF
2N8Jz0jvg4dB0v5fpqCWPOIkWpk/jKbY/AqONzItWuMm0wBxPRtZTTb+uXUjv2Su65029IanFj3o
x7XL7zndUkjTCT14DCKjQPdu+eyFCzIEIltu0ftrB1lw/KmPkZMyMve6eUIEHpBxM6WBJEm0fkN1
bE6oEllca8NxNiPlzztT7u4QT2HyZns8Y+I+o4KdTcA/Io2VBVdMWGMyTVzV+G9y91fi73TvlPjh
hO6zsfTEdVQTRYJRD1hgBvl7qhik2+ZTyDOHAzApf5ib/50PhmZGlEGCYlfWVBfjGZ0xAPpPnlhk
isWiVL+g+qJXYggD5oq381h2ZMXTyvr9b+SEOjJptBq5cYCUC69pRS7XTqkwz0AJ1oUlfBMZmvBQ
Ia7HxcI9dEW4BieW4VHW7SRkmEwVRxmF8LHMJvaWv+9Fju3lkPhgOgtNUqkxNmB9rDVis8LBfF6J
PSIczk9omjt3rVvGnZrF6iYboQKh/VWEmeojbmzHFP4VWCtkUEMmmVIKcYWOrvGV0Zmg+yLf4YG6
9+1yuafx9ANHajCwtIXfKufZjIe1j2yCuwGV4MPJRdBHF7su99ZexSx2qiq+gXHCCzGkGl1DA/3n
xYdM5ClyvjW3LtOC/2UNFVnFkeUGUML2qB+ppleg1/UXA2Gc6/h+5gfWxl1y5oUnqGmWEhx6juZf
v/A4bSHqZseT/Hl4YuVRoL97OcJ5wszydrSJPfuRjZ4oyh1oqIWQ1BywLaXvbUO7IvMqjsZLrfSU
a+8Is/ZbkUbYEum8PNSjiu4IV9ertXDMJk9xJvb02lNtWmfixYxoKBBcBFav73GAWP8IPlD8JfR9
8qJ/2n18FfFCDSav1Cw0N/mFZGP7gg4EDZBsT32tGDTjGMCLktTNNW3gVR2BMQWkM3sMxntoz42F
aDoAbusxDV1bqvAumxY1gRtbilBvLQeogxQDT0iR9zLi5Qdm6kLdIneuze9KGG6rcvtlGNngMvcY
47htsVhxBURKybLS8EE22//2ko1SXFFTMUu5zFKCzAi4UC4rJjkrFlLT79aYYSMPtpjFQs3q5HhZ
+d/RnGGgsQmHHXTOx7dj291wE0ms6cUez634KnyJ//e26nbtLSsG9cBb5r5piLnh1ll3FEP/ASzL
+BrznMvfhIDPvsDzE6WKyeq00Z2UBT4xT0EhMtCo4gd4U83JWnjRF0ukikY8nLzeOUixy1qiTEOF
R52oH6Vw4c+FQvNRmdMBKuKFz/vtYMZE8ogrgZRjhcLGE7BVjr8eDMLwgroqttP57+Aw9wlD5gia
7vHLSp2WZIa07zX5quRUjzH21QXZDWCnl1v28deBXgzBbVGz/w7H0E2ktTMv+NriQkU2Rz8Cfbtj
+ImquedKRezVyVPklgv9/rOGEAuCOYPwpBdBKghHmkW5K3X6S8n2tvuR7d/QIDIR0sbX88cZfZ8f
GVx5pPeDyHzFA+BIAX1aUbu2iSYxtxdS3su18zwDFP8y5GcoO31xzpq0cCe9GpVU1ciAktR0R4SE
qDZ+kg//DewscqqlGO1/kI3sPNhExOhY/Nih4/Q2U8Hi0PHTgSHko0rFDoNHuaz16G+X532D69MN
KeKSVu0cCa3j5bREWv/vG8K1Wv3l2JoAtAFwPn8n8F5okdHO1/H78NFi/tefRC1KdemAFZtWbruJ
c5H8Bf78dZFXMvqugaOUEeE7y1+pzn8tsLbOMDkIwakRu3SqFPoGDNOarNhFmHvqggAq8vNhSFPQ
hbsYKLMIBKbsRiwqtl5puO9USQ7956ZYHmCjYQOzBKt1ECplZ6T1TMD9JpTEHmjDUORu5DitaYgk
lYazGX9c4iWrRfiK13OiNMYMKa+/1FHnsL39i1wntVM/iVVYHmPVJBn5XPGhb23mW9+KqQ6Z4Gfc
WDEq6bSOPH8GoQYt0wUBov2mzEPgppHsRGOdRAn5f8MIKGt7i6JBcLk2VbzMmbypjzXpFYPMBj4y
UaBRas4iFkxKR9ecdYIB2YgdTSoDRkO/qPKCHtR9ovL28UiPjWEi2AEIqmHonNehsxVQSwtZKaWM
mYD25BoNQASBva7Ik0dlKc/890sTtJ5DBGLiL7iJAmbhK+jxIN7nnkoTHbFIzQAo+08hr0B5FCVF
jspNACid/n5uUPcjYTocinuiC2cIEsHxHfvrgqfp+4f9TpzggmY6q38d6OJut6QM5GokoQEnMJx9
3nSI3WGUlsvu7v5mywQ5+VNS7mBLcwvpcIDxGToXdC2ZrqVPH26X5SoStoPboF6dBZBmCF63++uv
ujwkKSF3SsFyEiciALZUSp+LLKevu17R+RHxdd1FYseLOGIx2ai/Y57vtHwoS2/kWn3YmyH8TWJQ
bW+LL9VxbiYSA1qIc5Se5JwcvKua20clgzuBnQh8XDv0Y3O7kYSmVdGikSFS2vgqQLEOmeVvGRYB
H8LdSiolJ3NckX+VDmSUms7IEjYoLuT2kNyFHzZuJGWgjfsVt1ZsmKQwujeHlBBdyt9BgSrdhqhq
xWPcBhMzwImy2n70NIM4vmcdRnPQMQcl3zQKBmfdm7k0+d3mvZmq+mXocddfNCYzv/itHsCfyi64
ARh9IXErL4/qavR9NiaILPHq526DZUlisT3NqdknojipqXJibHbJEMGVNJx8mnALEpTw9/47YSdr
rbwTeGg6d4tV2LEfZ+jqVTzD9sJkIxbrpDIWypXW0oOg3rT/pGyL/RggOqRy2GDh4AwzQVf1Txmj
OiOO7ZQ0aPtphnG5WzDw/WMF5JBET43x4s1+5nXvlVWLG8XNqUm/EZceMRypqHex57UFqrts1pGy
mva/oWbRQlQSDalX+owBkLYCuzkJnMl+JERhcWwaOynSQa7odwOh0T1V+RZbv54UIybkrKBytpBc
Ntw/P3/9QLO3gK1ES9ekkULAgeevR3koQHgSslF/2Tcd8+ln16twKGQ2eOIxO0PxlQRcPIU2lMPt
vdHKlnfTHKFmPkXqa7PVof0/pw/S2rj4mkSZCeYygCfhxrhaZ+UQkdra6HocXiWwDk3JfTjw0Eu0
CEbx9+0ZKQihH7zl93WEJ6rwNI7M+v8xuSWpLCcgSr3ulsUi9z10RuqqfpEwMiAe7aSlP+vNJcqG
qZbaEELVMV/Ibot/qLpzJvfsg6AKUcBJk2Ul2RNGtf29U4SWHZBBbwvqrD51BddYX/gEXGXLxsM8
WCdDsV/c6tsH6IH32eCWQI6ULPdAZE/EWmHCy8ufrfD75r6l7p9N/hGO8fXkvrxDMPTI28vKRBq+
0kcXYIIOAdKsOfx/mB5YGVf7zYBCSIwC7iTLECGL/OoXLbisjfnxrtdPew77Sd6geF0Ba1xuRFiA
sTN09v4d7540WsJ5jbkcttfcsJ9AXUm+IP8ZF3TarWtJexJJLxVc5Na7QRVZhNp1ibINvvfocgT1
AWmQK0ZCJN7UTL5E8fCzNeaz9MhSvV3lbZI7PEQqEK4gVCzEMm5+qcSzq6i8t2JsUuYluqJdi+pN
+02lSQfXhvxL2vhml7Co7hWWacttNC4Q+FhR2yWOEBDhia9jX9SBOefqS1L896OJKBiAsUADZyfN
EaPBsxlVGT5AWtgsFU7bFm53vU17ebu3jkgV/dRd1MiwjZxTGLCzanf4F4jSoaxH4pQQwMPlNGnk
6ekPjLj8tSs++TDXdDH+xWnAkoz0qwRR48dcpQkWofxbDZjR+vieXGlhAUCxC6th3YXYDb/7HUym
gl8EKC+0C+7P7D9aqrg/u7MBbZM7kXy3JGeeabBBkKZiYy9XBOX+Ih0wdVJLfcklFykSHnHA0rig
cJdxR3/HV/R+xmGc/eBa06vKLdmT1cErThugnPxRcX4VwOrdyIen3CjLycC955eP+hxuU6hmh+V5
FM5n8w0eccPk0gVwIdOu0FomdH3gRbCzMFDjOn4CJuWsX1v1bjb0k0OQC/sPZlkZE2Okynwvw8DJ
GDuj5GKTnu7JRJmMSRHUDG6X1yIuwZ4ssC68W5nHXs1fI7GRHhANfHQwd2oDwYJys8nJYYJc1FU+
lKKxaSjCJ9jVDhCpb1ndGbn8tnOIxrxeizF57D7VTI/tpfuuXXmsqNb1JjRtVCez3fu5rQ79WHSA
YbKOjt4ZiZu/4N/jNsR5YRydez5K53NYLOi9pDlZfybaJIJC8QCK/XqzKPK5sej07S5kSIvvtRb0
8b85LqY8wqBzcJVCkAjJhhNzi5qQQBPOvVNEBl3Jti8GGUTzDRjb2QxuFvKm7WzVh/DPuxqGw5Xo
vXCbfWSXraIfguP40wscuztKw9EkdTsqZz+IwFYTzcItP2B5DUwwoopbo+Wj+lmdNqap38b2bL2L
vqU/A8YM73il0kT2IKzbstbCmONlz1WT7AOBI4mYf6NGP+W8k4eOI1NZfKN8/twO3qw4U+kws13s
tfLyA/Jr3pwqp7cAcPfWmArFvkZIACdkaxPAuz6F6dxfxuN2nw+PGHGndTw7V2Gr+s5eQ9QZhucg
fLHl24q41EL1bvdmjxjGbG8UQjEuym1kfzJrDa1f1FA86n42C4DkbdQCuxKB7d8Ro18tUdG1qQVM
sJ8XtSBx5zNBdI1taRsvnQP11w3gTvT6jDWYp/ojDkhuNSdq8cIdS4c68FsXuMELgvVhR5I3f+D9
X5cymzezuHAVqh+ZMKLAGhOQyWr/BtOPyJ0qtuLrwmtqjr+epNm1eYESROyNmkp+K6vh+xXS8QQ+
KBIz6IdEB97myU2GPRynSY0h8d39XBdadLYkkMMBFOEUwiZDNcC33fGKa3475LaV4DU9S24ybx/H
QME0YeVOLVh1KXQF36nDIIuIW8Ni9l358bnvqepJXYRZAJF/g0+fMABvdH8WOgX7Y3SUZ+ENPWWx
zB2NH48M0QVRi4GvAdonP29hNN10HvthFxQewkp5KE9opGefHmyyXD6sAzrJQcQVgZa8PrNJAsAJ
IWfsqPUvKr/pS8YCbNCdBepM84M+m4MksXgKTidZpUvp7cW1oR+uQ9cPj+2ec/Ex7rtwc5EWkXsk
/f0Eagi4+2haiug4Xal0/5NtYkjhCVDI63NCob+/YnU4ufr+Z6OXYu9Ct+9LGoQkfleWDHIVTko6
bWEPQvv2CQqTfecAysDsrgjmY/K7aUISumLUPOW2Jw48A8IWr/mbMYSo3tvRjikqLawLrsQBt0mZ
peA0pTAJ3f/GyhQC9WjvlC9B0RC5TrJ8IU8jgUDjU4HdIUleMnkGnm0PD98mJFRLnVLgG79ZeGJf
1dD4CDRy8nmhyPqeUknsAt7+I33Hthx63dnGlZH/jiQYQ+EegqFDhZjCYH4At0PtdS+e+ArWk7LX
6iDozdPEBAaQ8YD10hs2Hq0sca3h6rclfPgvRDVK5Bq0VehsO3dtnZGRzJ3Wr0sMrNTRWog7D3kl
FnZ5T1fOFNsGhgMCJrx/jg8WMfxEq0SfDT8hO7LaDn2ibBkIN1DAwuCIUNPuHrZXEaUgHJrgmjXU
SJEgDu8S4I2g3CYD7P91f19dqOBIQEFdT14nUvBGZBIc200FsUzz9a1SMG/vOW7/R3OzGOtwmiXf
cjVe/DpVGf4idw/QA8LYiTQLVL/ijTwptg+pcFsmjhizPeDaCga5eqex0c0lJqFPfnOjEJMjd64b
UiKcu4fcl/rWtFzxxEHnWQ+AtBeP2w4yamL4VS40giMhg5liTxOwlcopyAPLoMOahNWqBdkVT4sV
ER82qjZMkZtY30tvAOjjd1I9HHq1btYoB82DQgz+SfF3oTm1B6DFcAqNhiGkPoquWCHPPYmXhkeF
wC/x78P7ijtHS0nN+/Cu9MkwKCdGCgIj9NruuOrl+GmvK1Es7SSU25RHvBIBXQagmqCl2XCIeXLU
qZb+m9xuPGF/eLZ2X7VBJyCwUL0EJEg6IxyWdlDFHNi+/vpTpM+S2J6SZgVvcZ70/PlP7DbtWbn5
+nq1GEieTB9AWGtdS76luTNAugOU0/rhd4IVOH8yznH+jW9sp51XG/p2RCoSZ2CGjffXWBxcZsqJ
JAJXFqGVCGjRkcraPdtHE2HzvVLG1unFPOVFoQYDWxTBN07UsiJBNvaEDP+6q9ttyiEZrPy06xqo
nJw4jLgphHNfSvRp1x7vVS7pVpMuZ2euwQkQ2I/G/EUkV0N2y9Ec1LXP+y4ggPn3ngDz2hpiuTe9
ae+bnYagz4YcnyPfbcG9OpFNU50H1sKlwQCoQ2ycF4uBSdQTttt+5xBfEaYJlx3dnADURJQaUTH3
zo5A0Xc+cDRjGObDtVloJUr2NtW8862jiMmeB8lrVRXLoTG0JeLyHFMpSE5QYPsmLUjmnDu60sIU
64d3XHNIk198CbStduP5oyALp1epP7WW4Yb1iF0L10Aphma4OTq/UlKVoqu31xJoTr0MxPWY3Huw
0tdlbakucyimEseuYlAPEXbF2p18gOBPOcr36+EcsNRBVejgzmaXKGSERBP3IAdHfd3XGQOJbfhV
FBYsvZZn/k+iKA+50TKG8Qd59mPNSQbABKmkXEvqZhins5VqwMo78Zi9MbbLElueqT4Zba26IrlR
nofdDiWFVPB05UchmtJqyljmWq1+LUuryqaRphnvkjFTZxhvTILIauadp8VCboE/eMURT/IX0z/4
IQuiasSePkSikmw/NZ/EkYtHBxJYzcwR5ry0gOkAy3YGlDhZlDIWkKlzovbkwmZboASS1ARFZ79d
oZlZZ10q0trB623ZP/PPWf8LfY7og0VPr/DAnJ/OY7QvKUbHiiQZIjhRuRW9GFA0tcUGl2K4VGSo
9YW/A7w0q+vypvQgiI407csyPlSorqikXbLc5sYAJuP5PizAL+EV7hzikRoGjIlFJDXgNwEsfjWJ
OBDF2iwotsBMin/ToDAtJii6TDfie/NJ8TTUmRcmMjhOi7RSqMOzw/2vNXmZx0tiM4qDNNqnAL0R
/QdrsPSYJdQ7Vt/yltR0Uk3yxvZOp/25SsyXHBa5B6LvjLtLnamGP5bwK3iOKhQVtaho4CLcIDcL
yY4CAM10c2+hioAIqYjRmDA+iTE/eBXlHDwPPkp/JUYl1uMkvmO3+vEGaXzFX6dNPWfclY6/+Ttm
70PXJgAnXs26qMi+BcrAjboS6jY2Stuz/bbi+/zCnzOQ3fH6sDuzn4n/exHzfJ/duIUc4R0zEOkq
R+vhRT85b8L8gLMYPSCMEI12cruYymUD1HXfHsjVgqN0OwdVh24xyNYET9Vx5y98iQkaHQRpwiJy
OWXXinePbZ2MggHjP2u8EvA/Jn8q4SNtgJlVHTlJ/Nuxa3XffxPbW4SJe0PYhCfrlsjwMokh6sE4
s9IQ/BWrsjPLyScz8C1VNk2OFsokVEbUlNfRfGrwbPByaRD7CThrRveyHpm600NgKod6gDZoyjSr
OaUSYqeM53s4BoAnIK4SMHZ3v53IN52yxXM/ecYQoe4v3c7+XHIqVE+1E+EDboGKsQyuhw3lzR7H
v7CsA6fjRsddjSRIozXhzpmVDhgg9xXzhZzJ/Gyu/iDykdlH7o0UOrY9scn4YQuT9UQPYulQTyP0
+d85MSObtRjXTt1jKxUUyT4bEijHlsGR2+avuxO32O7Xwi2ysrbJiZTqGnHckLFnCvSyvf0pjWWh
RZ6jXVW52GQqAGLj8mgX4eOrRz0+lTLal4CEa0fY+29cTM6R8RErygOtbfdORdEcBcyq8V5OOmHa
VxHpo03Hb65vUkyjqwj+uOsl5VMGUM9n56GK/llxEjTQ4nmlZt/tPbFIOk9cUOLwsUYgVOnydCBh
nFptOvAlq//Z9/cGJjc0kvfIpMHFMnCwrAML6598Dy2NXV/T9vBP8HMI7Nt7u+7rtIlrqCsquXe9
YfQZlGqtkVrIztVJm7NJDo4Q/5cnPSZvhAeH3C1dhMJuqrCgR5GQJzhBuC2iUMYeurNtXUAptJuU
rqi7hPSZJJgGn8yeCkPk+clKx25h7nzWoByoaP9UVj7srU+v6qFIRaHFyJuFNQQF4Vkmr5rfou9s
DGqt3RZTIPHF35+O4Os/OjRf8c08DTsIPnoKNPtpIWjrJHR+5IwVxg3294qB/wvrpfwda7ARCJtU
CgTWHMU9oEScAZGiYk6UO2rJ9J0F5HE2HGypE2IQqVQ8e8fErKj/CgMJmQtCNVzQs3vC+RrbqS8J
0fXYDRZ4abmbthdmb0dYciy/cBLbdMP5qDEm/XmdJ/EhxWEdfMXryZyleSXQEr+kS2hIhIxhVHkk
8SEDjvbsDPuC4lrdQdgavn3Ka+JVaaCsGdNalv6nC0hGxpmiPVBNMuMGK9GCjKBXtM5C3XXJr+IE
lq9WX+yKJ3jkTFS/HwO5E0NRnUsSvSG0MaynjQnLETAsqOB2SquLH5WTIAeSsOde3UcC4g4nPGnV
vzDVevjeCTbt0Lfrnmbq9XZlJbquKUJv18KhqsqbK+cknhCD9ZrwFXMSt7FqI1v2Vqpjm3YdMCIZ
3QNbOH6qtYiRgp/V4F7odzuft3Td5aGzWz0HKEGwgPOpOE8KdMxrVHT+gTElc2P5MVuEX+nZbpi9
LCAXQHxVepwYWoVVbe3vyyU/7u3ynL3nzjQfnf9Q6a1K4bNM9u4NHUE0MygEOHjP286kjK69mbeR
F5Ps1Vitl/HXxp0cw46qHqpL+nD6i/aV5XZjHXeo9pz4KzPuJd67oorJz82sop6uvhALezStp5L8
P5FvauMZ9wDXRDFP1TLdwvqm6BQT33JtHunTQy6aDjyAIbN3A19LDvsc9eNkyNLc3QXzZDiq94tD
4OXFcOktE/wv7Tu5ATKAqs/p/QZu59RdZ109XCoczKp3kuqi4Uf6UMx9FeVDMrcrKKmepYy2/s4f
f7IUwfn1yQSyfYx2oDNPKNqyXXINiojfcmNqXhZRfWFxnQvnHsIp0PwTfYfVGdMJoUlG97Jz5CLG
HvUaXqI5pymH/th30Qu0X0SUlPgMiTFSqmADLo/NKiErggKE6Eex9czCWJ4vzXW/9dnQuHkRdysu
bIV2vgFmKNZWcb4B0FI8S477oQ7o2pLZjO+CI2dMFskc56EfHA6KgTPgiQam99h9qCXBNagogOGk
pDXkC6VUinlKSefyaclvfodgmPYuJj5UB935APT4zdX3Er/WzIrPM8hOYKyrYyxDwL3OExuPN6UZ
AFdRW1qf8l9qtQZym/2kFO7b1TnFP2pmguuGPnTZatclxfFR0lsigVe1bIUbQuL+TGNHf1jaKgHy
PsiBLGz3P5KSdjDw8UHST/1Pephm718HWjkQGH1s32ULTbb99bUP8wtpNVhjqD5NyZYH/42PHAzv
eFNdbxIdPHwZkRCoNzOESBe1ZzQEH8zjuUsfqhibUMPJ8OTcxVzcbMgCPuUnIKSJ/+SBK/j1QgBc
G9flKqm/fmt6LuUp5V9U4JPTyAD6RO118vMioYz1PGn7fNac0LO3sBXefSRA6d0qJ50mu/rd9TTl
XzZpwDviZr5WVj9zzhuey2LlukUKt1ZEs1Cpp+eXj0pWdnCzPuXR5f/uTVohi94dOATTFRHffRry
BhHh50p5XX/7ETI9tSWcpmA7U1A1Y7BDbG+HESOCFtmXpyGgRXe55RHljpgw+M3Ryl99XJZsJ5V7
9rJ0AVVtlIohnZEhgcUka64/uM9oc5YAkmVutaM4tCC4AmTp6jey5WhsTcOteO6z2STdKmZtFR+S
YTLUyfhoLxaq/zMoENH7eq1Z7dU/QSuUH0JJ/3aMFlOI8INGtZmkVi25a1HPjU8bUqn0BEZSr0hJ
gJ6fyqUsEg9l/+DwTwl38hmY2+IO7hIEqqnfT/f7Okoarb8KdY0o1RCyrOoy0Urpkd7MM8HCSa7w
puX4iph0gyf32vroHdlEiKxyYfLCYAH9KD6CUlM4CjPivnrI/5YPISD5H78hTvxId6cclIA7Cx2Z
RkA0OEBx/fTwyw6WW42WcnPwTi3nOTyLBKF3M/xlI/FVYpOa5MiusDd03GGcax3xI2E9ERhKSGgv
6S4w4ZsSge3A95BD2vCRtAp6w/SR2DN6SRyuaRwejvaZKi6U2EmQjEoXIRvGhy2LoIJecZ2tpymV
I/cMJ4R8fE00HLpt7ZmdiKwklX9taoPbvG4rodttlvBp+9ak66T/Q022nqNi4KgMQILjKSXN+1xB
hfLtd1fF+G4EcB3OpZxDkfCtg+BZH7YSOUd417aD1lg9AXo6eMzXtw3yG0WGBX7175I6GsxJdLD6
Ht+VO+JMNT2tqTHFH6+/zuUaABYys52yfAG5yTEpYYFx4KfhnbXZ+RfbZofIlxlwpFrkmrSAzfGF
L7Ibo41jZVQ3BLaHl0tN67Mymmj0XsE29fCWL1GmtEih75MOShUoD6KFSner/hWC9hpFH8pIXcyO
3Flvb/VrUpavvpJ1sQjvTebeGQOg92wr/yCIaQ95TMev5w1XjNCgh0kFNtK3Vaah9Ckq2XB01Ia6
7xt9HHai+8d71D5YKpzS0BN6+y5quRBjWwNS6CtY9Pp3JQj5TUnpUBjaXiibxFxeKx70eBkwp7nn
oNZUStUo8M2CT3VFbXJr1hP4AAHGGS7a7yW5FAkmaFzghsXRzEdWwnv3vC9ULbRudZ7vQqQqj82o
/2cxZgalixqBSiCXXMiN2RBBkLWCJYnqdfcsf2kk6PJ7Ld3CGaZ3TuWH1BXxY1F1PoYa0jmY8ClX
WYi5kfbkRe439HJb0lhY4HsWFNX3jefbnnt5Bm2Yq1jIyoY+qaNdDx2a00QN5plfJCPT6moM9NCg
pMJ6ySDVEjtpl9mwVhlfEIsS4NtPOfaJHsAM1tKfT5qKTzqyBGzh9OI6C2FRYklm2aDOFi03S2k8
b45p9pnDLwHBnDZngkIJnNkrtSsZQQg/wcD8PIQIvVuGkUEgmiwzC0CPOLYEtySLY3uJYxOsCZIQ
eKr1d6vNACgJYDY3MGeBlE4CIHpUd/9yJwoUWpKoWeAkpOt/ftIsmqMGLQhQKtBx63jk+VjDXdKs
rcAn3u08aSkSveh/CXvPOvbF9diiT4wMZHtBSQAACID3dFdlVa5B+rdk8tdbhbERREH/SPpquYUQ
gtCYm3G6tXSYYnHUnWLC5qLwqiYzfvlqCZT8hrUGS9PcoCsGig+BuwwwKzIFaGQycM1IvJEKVwer
YlCq9ljBqJqUspDjbdsAPgv/g11vd4j6p8BgcIKj8kqYumOUZx/M4oI6QypkyavmwUdSZZiv2fzL
PHCKCDlGLuI7RKHs9Sk2cJOWCE/nKu+nLCpBTG0lgxrfXxujPRn+MG7pI7wzRtpaeayUysGEUKLG
DD18dsEEgYEIW9/5m0In3VSkoyXwLnUIt99FMz32hRetHbwnWqRp0BneT+avPrZICOBUwQqN4sRi
jRYU8S64UZo5ZEvoAwTv/54svO0fx3MyXHAkQj+JY9xSlqSTL/0MfcBfNmdzhN495cNt5q0R4fBi
YoJWXzbFQpPc7PrFNzBoicLJTzVTwLvK1gaGAgJ3SR2AOgKKnlIBdE0qZsZaT71/IWGo8TmEmyyN
YJ3R3gdR0S+bxwUhv3gbqBcSSky/MFJXqvEtlTGu3G9pr1svlsMwzKiQiSSC2DOiOdAVsrO8q8Of
yrDdL5HaGcnyPEY+Uj54y6aHSRmjSirXCNil6UUwROw9gyNrrb1BWhm6t9TxTjpqhAouqO39cVox
Vu+mVmavpOBFSmysvwgkBmtinltpNkTQnQKXxZBBBJRabaSRoB3/1MBLNCmyQQG3pQGIQcyB4nZb
B9NcXmczI9jyOAV7x9ZSLcCMQqlHdgtEINUOkoggQl1LM31oP/c8EuUBsCcSmBmOjnOBqXfCrmi3
ipghmCCyG14BKGLYwCCTC7r8qBpiQP3+Kx0Ul5+6KK26PlpwzRJyV208bzDFUe86222+ijmjleX+
xVi1V80bDNrSx8hMfolUKt7s7IdoAKYIWIlsOjEqzNunYWmsVeQMr68yasKmlGGRHlkkriNeGoa2
bkW9Wwx1toazH62E3et2guG1YuKQIXrd2994sisCqR1y30+LTlTMPcvt49ajTcde2CeAFiwo8jjK
NfRqzlnEdIJEfedaxZnU3Jc7nBIJ97vOJ/FjyQNpXHuEJaeyPPPrgXj0ljLCt4TkoOS5d4mF458I
3cCNrz2h3wS//AuNfX26CKZR3XC319S0ehfUT2rbZpBHLVC0wturnnbf6jqNdNcY8ET8mrIqS0+l
xZHt6BU+30iuiknmWamUdFkHkGf0socYGiUIgocJhmjUxjKT6zHGIWHRlrB1x4lgjpdqVxaGcFkE
ZQkANrPh7PR1e73ees7903ccQbDLk5D2ZaUxZ8bOITlP20a7tGpv+v3WVqdEcQKp+fMGf/odh2Km
ccuIcKCNr2EW181xBWnwFTKlDVJSxglvUWZXQSk7AXr6iZL9HzcNDxm3hAnK/OveUC/ZdEHVbpKh
cq2oXKcGbRIXmLZMLk8zJRv2YYdC7rRFSzRD3p5bnbSLFvnta1UCNQ2DSTjxaI/Qo9K8W6b2EN7B
lSGVMBGRrouhjsSacnybjLFWR7OmWjywhrZ0fIVbg46qMeHhsiYVjHlsOFv3dlkgS9RpR3OgRS1q
+ZwrB+pYsdQ7iHWATciX0jspXOuuwrzWnrLB2viHRIRj6gT79HhfxpEVH7v9JypAPcqf6HB7OJFc
cCRlaDBual2V2D9GolQapcK6nuSA2pCDzSPiWbpXr5XulCjr/21eMzpUkeK9YIqC5Va+K2j0FnXI
B2srf/x9HcCxy6E616LUPcLx3KgdNYaI4TyFCpdN6l/bh/fNbm15wLXtH0+t/prs1nao2bDaC7zc
oS11iwXe291IFjfa85rQuLUQTGeREwrpzR0Y9Dq5F9YV37ZFtigaHUgyT9NxmsNad33SnvQDEEBC
R2ledF12bvEaQqwbSYgy0nC6Pig0nYTNqIAfIndIWLEefGZjhQ9tRJB+wOYSropJLOyIQsP4B33t
+iIvInFD2pnDlB16ozvjS70HOa7TLjUgA+vl0wqjt9FCEUOCFmEghKFrZdEBpaO2nWed/ZYUSHR/
t9rTLx8B3ugULABwm6L20DNj3Vbzqam3YlMl4+8lI8W+NB+9srFPjHjFrjbKWC2n28pwefLnb2aq
kDmNk8IpISdOSdPMWcIPSINJgjAJ3vheZsHMWDvOVfrbNCnaUNiOCC6XlMaZEyKqJt+kimtg4okg
BO4iLdXdX2SLp8ZUbuYAQhaqSlIaW6zvE7GbZn9sMdsq5Kh/SOr46t+vE6KuKlnCeilJF25HpaI3
grikvQ3qWRgDyTGROcKNifgcPczxuNNFf2KKSAor/Itx8inNH59s1KJKzM6pX9ck0GmPkiG7gfGv
avT8+cy4nHMbBmIBVLUcgjNBcBNGVOy1H7n6m7vxlYrGmuc16R3IbVYgAcgQEGkgifqqEDC/jcdD
71Swb9y0oj0dQcTy+A2EwqyZuMlxnLKO6xQ/8p5VSfJYYvYPHTQk6eymxahrS442nd9WbY2U1n2F
LOCXjSQsiyITGiFgnlZx7MyUNk9lYtUmkFBNcEG0odzp34WNG+Zn7pIXSfCo4pbQozvN7TUHtxJj
egc/EW3I7MzxQI09Oo1gtHWHlolXM1tL3FULq+9rBUw08OojzucN7ZkyaX09XZBzjJkxUXkQPDt8
WgybNZ74MQEs96PKhdhaoxmhgJab+Y2megWGmhRZnWE7hJuUPmyHtJV9xGD423jKmp2VLysTPjsg
o1DtfwrX6L3wsxxIAMvfpiIxi+3XazWWyFXId4Vg2qxNRdw6pGvWOBsTsYFy/HTOsqRL/29EP8ED
iX8mdQFXskLnX4kzBuJm2RE/vW+rYetzfgNPQ2+roXfQoPmIMlDVxRtrPqyqZIUCsDbzmBL+GYhv
OmmfI8ak0nHemmYhboNVXziaLJ06tgS4PiGcC5pecf9gTleL2WeRGdieuJ7Y2061eIQaKDq+HJLp
fPBAJdBh7lKdH+asldZinGXgkGObBXir4URkafS4d3f/ulAPOI5SV5z3Oqh4EH2HUgjDXXBTvDY/
7Dv0Bl+LtxnDVcZZUVnh4h7DruZAFYoDEt090DHCpdR51mR8PN7alcRnULPAw9Wn5YH37Yuw76oM
3tuyrxpwmV/o2C65kkbptQk8uH3sZV9S4Rkj+6T9wF9ENlf3KmN6A4bWLzx6NQRmgGKLbpyAH+lr
TRXyEeHaKP7mhdKyCBK5pSZdlFlnr7jFOLebtwSZlzCxkLsy7VOS7PEzRz+Jw1rToIrJLRxkd/qN
qbl5raXAWLs8yP8TBKglzfZUBHhC4fdCGPIpSOZpXTjNo6xmyVqyR53JtvAstv2Q2Fv7wtWDJspn
oZ+MAFB1F/ZcspI1rdRwerL+RReMmrQC8ezb+Btzjihvu7gfMc5mupIgZGNIWQeqsAI8CYyomL2O
xEVgroguEGo7E1zoyra25VqLaebLzL2Te0kXz4JfRzEqswRkXHlth1tIJNhJDXIhmtnrTTj8vZgt
n0ykIaiNo3w1f8QNTtHtNmJKcDxNCaUO2OZ3vnyJuY5Vf46PSch33FMXaK+ffm6/g8VUTWtl+Adk
Lg0oPvH1NVIBn5TIx3XjJ4iugLyymtEb6xeXpkRmU39AOiXdUaegKuhc3hXKRkBvv7LQAJWiXRfK
k+BXso6An5L0BPsGT1nckxh+ma1vrFpMdnQF847VLimWsdqVaRPSxGZRJ9i1F+ntZ75+AE4An+3L
kbx660pZuP93E3nxXBt7PphkO+R6h3v55y6MBfU5vE26OWHpxtNUx4sOHxnoPO5Zm3Jf9U3yFWNa
/u9l255OiC0re6YrN21E8KystEQ760GMwvjO2v2NzepEffp47NK9r5MgqjMEZtzq0idEA2EnI49s
kQue3HRAoSuiUYDiSoBRL00z6RXu6aoazgQBj4rzDwWesDXyik6mL5/oMu+ptDVMNnhRqR5iyhh0
ZBKLiQbYH2BOg1bOPW9u5R4te/Q6Gw6nwfBaKvXY2NfIf7MxO6ltDNU972wGMSD2fGxTlkKJeeLb
271wL3o/HEBBov2DXvjenERig/iefE5f+eaPQMvCed2bQGOOd7ApxoxqIx9CpGlEykNoLVGygB87
jG73tmgC7LLbIquPJ/CyhCTSdkksjfIFtTunNanhahEgWIC4XxeA4wZ9wRcdKqY26FNbckRuzv+t
/5UN5FB2XsMW3FtR8BFwsZkBMESDTv/jv8ShphYEHV5U1p708qLv9Fk11fAmu8Shexwiod/tzRUj
NP4wEeJhIEc1ZELx/snj9uNkd/h1CZlTYUmt9OHqvuZ974Vgg/4lwQR8sbObus6Z1xUkJutd8VuS
nVQynocW+wAYvbWpeOoJfDe/U0TOEkbUcQRR2kj3PQoKZ6ZXfxSbPaE1qqzPRZRK0JnCHzANNRTd
0VnBxtrjtVuzz6BQ/uoE0cjxinUFj+aEXNiJaLBZciUZjg+DA7HciKchX2LofsmGnDEQ21XY2MQy
utt4E910j4ygzf8S9H4AZ4JHN4HDQN0u7uBgHuDBMHqHTQDXOEk4J+kznP+zlH2B1V+zis42X/e7
+/pJ2BGtbZZZvV3hkhJKo2zNyT9Mb28Qz6lmw0ljgK8YSbGqCrAoC2jK1XQnrDq2/B4mfwbRh3C/
5N0Y03RZweOvryhbSoeqcautM1NWCYyJNE05iH6oTU3xFpYXYL7t9If+SySarpYlglO975AWA8N+
ijLxkCvsrFEnyuxA4tbhS2BtuE7bUxi/PPEWRdS7tyr72+x07DmBY/qbxRo4ckl2NaZWHVXxpiBE
PZVpofkTebzLgRhM8czCCzMhlKmDiwJ9b12Wuy8aJioh/ZcxU6E4Rb29ZVd3c6Q3Dn+mPf325B8N
Sf1zEVuEcu/ER9QbQxV+wB0o8qs/Tj16+GTDbQNUE91kJjFX07CsQKKiWEoei+ADbV8d4eIvBOBQ
xZjDEfkrjwlQYrG99lGH0gGy3iq4RrIcO0lNrsFgVMUV2J41LdydEqf9RD4W2jgabZrMtiCPTQib
epI8tE2sMjKVhF3eNbj7Y8rgPcXNShA1HXo21w9ZBzJ+9SNYo22BEHEjImv1A+NUiVvc6D/KEVTI
A3qT7rDkDEVimhdliRjNJsQ4+o/TpbAtVtntuQHxIQhdnbwYQApZwVatSFMaTuxGuPICouMcaBKn
BayRuYzpa7+11TYRdXDX0eC+mPj6F44tvNZH4/ilDjE3dYcqm+cIQHGSOPR+GQw7kcnjd1DlZMg9
VCprH7Y9UPORvr1+K2wtbsKBVo1bJTrzBENq9bZLm8CCNyjCP/5KXQ2WYlLzQSSzE3wzTgqN31a6
1WH7YxE9bIK5pqqI7UcUtjJB0JdWPoY+B9jFSgPL7FSvAfDsNr9ugYZGe73rfAM1ZWuYbeDr7QR0
4ynAO7qGjvJd3Shgx4R3rAOhq4gRUfrOPK4DCnEPzftD1xOsheLWbs7j7Bt9DWftsIfV+u6fRJ/M
ipK64UIAYPpBaRLINLGwNoArT7kmFPaIzDrlAwoBAbSY2TXo1LjMiGz4CYR5G9MRqwquUtgpKlwT
RAn2kA7J3sX1rplWlDAWASVgHA6NJhOsTIg4EEFAHdVK5Z38sf6u80/IYV5m1b/qTIPGwCn4V9To
DfZz7ZBR5PGN9AAmQ6SGwFBdyBEvH+mBXw+eXx5CVk7m/790759tEiYxr/TDTI7d+X+RhOJpt8lt
rWUqRbX9lgS+gFqxdQpUUIXOW810BOA3hPzeGxPgWv5qQ0CC+0EWUdjHYNLOazVwfqTRMTGb1VvJ
81wQWbAImZGrvWqnzXij+M9iztBty2exlba5znYJeM+H7G9dscwFRZ9s/qy7hDU3Dhxpj/n15W++
ObGoJyj4d3vS4c5Au1SrN8+Y21eHG/hazLdKjcwEl/7sZLzymJPd8sFwOCFGMBJIgsk4Xsiszmtw
EAvlWmlc5Fnxe/h/gIenBElBp/ewaqtwMedDLArG7fLSrdfM/qL7luFERoTen8Jmu2PChf80P42w
ZgHw8iMsWUqZsla8umYGPRa2T+hiEArK3D5Y2n3s17dgcK5g4PLZRAhRNGvlLSUzjqs9pkKQm2C0
DDQdUY8BriYLnOw+gXFaQKUAkjplslJORwCHJikitobSeg/9UtuEaleNUVD7T9VM9Q/QPC/3XVP6
xF8hU1c6Wo06ugyTHgfJgsuu0NG4dmkGWUjTaKQNo4rdgQx1Up3qOhIvS5WC651ajKKyXehjR7Hc
D3hRBORxmd17kpnsgOKUhim7CO4uPfO9FQXVIQ+qIUm0Cw1gepGovxeJkVq145kvG8pjAIgu/i81
W+JP08Bfuox5faJz7dT7HV2b4XJeGzcLoqHEHLuUMns49bT5vpesBEuAROdGlcLq4QmAf8MrEhSx
YE++pIfsEE/tExCbb4dti9CGXrItDRWJ5gfhnglfEhLncATmVPn27Gtf6/siiJzc6ArJbskJz4LH
4UamdgHeTXkaLKlr4cv7wU8ITtzZaXCvVGXCG0kNgnZTanV5insyh5gl8Z3a9d0W3D4D542wW3Xc
ucldH8jZyIXv2tWRUWP8o9JSz5+HCwd8dyb/BoSAhK4MykUIQ/06JF6VFL1kzQuNHLasrsi4BbFa
+MUFHwzxnOpS8G6U9uWOnwB6lQraM/XDtXZyT+0pekpeNPYIbDk+eoIz+VAHrhduFVIeAsOqX5ZP
vRfumjwfza5ejyZBZt5aswVdceZwVVFryrJnIjPpYoUsMsgdRSLmUc3c/cAErfI0fokn4fwAM1RN
RtK2NcdhqWq3fg+jqqtn9JJmpo+IQkPajiB9iET0AE6HWnSIGKs4dMbY+VRr8KY0H9aoyb4BfJ0Q
ssx3bQn2w9a2oHHqqHGSTJc63nekZGWNF7VK8Wtpaie1lIG+KOgeI3zsNKi53502xkamUyKwSJYt
3VJUa/ZySd98UieAeL2wvNPfU5vQ46mGUHhOYWNI3GMWNck840cZmLXSRPsRr2rIoboesl/wg4V+
k9l++NBP1lE14CuvNzRLoiQruZwEwokisY/c8MVK/9JTTvt1wACVy+c7B1vYvUVjUieC7fsgwZ+Q
7MrKeh2leifcGabkHhBYDH/HD9DbaJWrZ9DIDtmnQ3lHRlo7nNKF3N+Nwe5GalI8x/UaqTbfq8Hk
E3LHkbICZ8tOGbe/CZc7fLoAx6o+y3bdHLwZJtvWOA1NTLTXfqnU9u6OvJib9CqKG+u1HNBB8Kg9
HMkOf6Y2OfwJEXcg2MxrXyLPmVmiXhJNy1XqNaze6j0SLm7/RVbpAiciY3Tn5+YS7jlAK0QbSs0a
E2ctn3o99b69iPiLvcXbWnI8NybBL5bkQzWsGv7hoq/S5iZCim4Jn8IHNwHR4scug4XxU1jp22Nh
zRBAuNSsRxS+J+iyhJgsW1lwdyn2OlLS3rRncTNLxpFCZdSlrupMlPeejqNTp1Ycw78vhvURTlOl
E/9Qo1mGoN4dVQQrlqw1qOcTH09u7HRGmsFS/8WHoNp+lV+QSkAURGxO433aPUGkQHnIyVbHh0LI
p1YN92FjDg04Fej0eJ/ADSfhYLVEmKJAz30UVNTweMTFlPQc1ddeRkQ1zMw0339Em7U4atdXQPli
gHGHUVsG+XYHWLVDCix4DiZYtXox0Fash2EWKc8/xlpGzbVZMNO3fjbqD2Lfrn/MiBzZtyEWzIzc
G/i7ckJXaADL7q2tDwnHX41RIrLTZxwGii2YRNb7BKe3buBlWBrR7Wfpg2RymAw0zi9bUbWSBLi5
q3a4hNI12de2LGhFoj29H8/pJwOEOnUIIpBHuMI44FzJ3RaFGIHu1usvnneihTNpSxmqtGxPnmiF
/NcBG7oDqB9r8XiqNMQdLPGdXXMHl9vJskGLQkYKdAZ0l9hdGJGbQAXHlbWgMEFWqFZGqushITpx
Xg9OnFNEHBIJX7I2quO0HGm2/co3uqrIJS1OwRimiQ3usq1nKj4BvnWefOSDKj0YafneJ1tfXH5/
B8VnZsm97WBiCr/6BOnX1yBcMEJmowgLo145xXojKQ5YTExPGINNlkt+Bkapx7D1o6J/m5itOAqR
wjtDxh3LV5LkiiuM20mcFC3qkfmyk1bMKA0kUQteT0KvNWGhydjudEIuLaUUkEZAUuxnoqV1t3dZ
QOqY8yKrlTz4Py99jDyQ0XBUD+QTrFhgMjH0MdDPIK+qQ8lLQJjJAJ16AO8AoW01bh0I6Sy3qIk0
limsDZEhXalbwJXr4EtC35dOqpAEg3j1zvsASc2H5o9jubKrNp5vLMMd7E7+vV/sK/lBh6Z9bfmT
dGbzy/PGQZsfyB6G3G/H0RmqeQ8h8P/exNddl9v6Zo7GHCVrpvLSDP3/FThOTX4A6NAMW5O7x/q7
PfQv6M67ULIVGBzjJc2VIeLb0vUtlqDCP+PSsjL6y3WtccnTwqe7uFpmB1CHGK6xOeS33BLQVq6T
dUMERrNRWOWZRqGrBaDT3KqsnERJk6OCnPUt2wKvOSxUiFhdkkwJ56uC+hwotOCTlcFfrgDb1Frg
RwWU/gH/SObNkRAQx/Xrgd1TGNaL+MU2I5tA3xg8YhLhWz4nBIBR/Zt1uBRmRQM5dFfsKdSA4LtM
XOdrzUjU3a3fRysj5ThU81jRF9q/bTGQcm0EbHwU1e2uNxXHaO9/8osbMnbB/9QwWg7VTRLoyFu1
EKGLDJMdT/HYpC9FgcKwc1LQOCrYbCeIM13iFydC77nml82uDOmQTTLq9kmoPDStNKvj6Np6FDpw
dhusDTgVmQewFkw7CRCyZUzaJ9xp0JcchDfx+Km78AofzoBTBQQpZgwimOfVwIvdhzzZ+vy1iq4p
67/W0HyAr3SOucDPZwIV8GJkeK0Wq23rxBx0+X4t+bLD4nFYcK6+8o1jJTaKuGR2LWbOsu7BOhPG
zpUcdmC4X7QF9hct1nl4KPgGs6O/8mPa85DPeWyODC3EZMG8z0pv3QXaZ4Qa2EA6KY1oDLHdeF0A
Lbk8QeH+tAi0Vj87DxwiVhAqpGRBAwzwEFGKkAe0jmVJjbTH+DuAOuSam0YYbaRCBZ23SdniBPEk
G3xhQy4pqxi3om/jaPxHvlOf5gUgM+TGnV/8RsDa/3u9v/O3Q4l0z/gKHnwIebKKGV2O/HxqsM/8
YHV5ZuIwzeJFIgu/Eio2wZMztCG9iI7ZJ72fU7h0hdwKxtVYm8KMKdW3dDxGKlI23nyWC0iE0nVm
5dM+fWCy4wcvlVulfkXtmuZBza3JevmeDwFEES2LH5Uy/16siO/DoIEBhfmbdSjfugy595odS4tf
ij+Kge8lNDy8mY4slyidjK1d4ssykcCR1rX66GogguXGCOYhH7Dx8kz3DeMa7CgAPQAEObbinhmL
czADcFPHUDi0SFTCq/Lz0dakmAh8hKtrZX0V8e5xKcu1xi8QT2ZmDpqUyKfQzoMi9uuyx+mF2oiJ
XE6Ial6e2BAVm+oSKJoNcBedZcRf7WUYm1HWrpEb7Koziw/5zkdFzX4NA5k+6coTJzhl28TFXggV
Ua4Rq6+aFbqPztL7+ud9F/ZnYAsD9zmDybcnN3RDxQK8JCctyGgg5BD1yeocly9LFnwdY2BEFM9e
QJnxCVABuW+ojKP1J8Yd4BE9G7xAjxKncxim2/+i06UUw+VN9rkhK+oAlNmhkgMjiZaqj2XfQ0qY
lkwok44gL65P4agnOwcihK6zZnW0S1+NVWFOki/lAIhGTIop0pdPiFF8KEMqQr0PfWWqMUx4Marn
jv97FlkriiuxiSkodNFbIRIRVIJsjOhOiZJQe4shXLPmUdzcQ4ZtF01quF9HcMKS3Kz4VVHYmGJY
L8l4+x16863c1ICLFviU8cMCWOZY6I33aMxk351W9qvpPIvJJI7FRPHbPfcj7+dpmchkE0HYlgSG
zwbFYdgBTyNSLND2oHU43GotZLqEVkR24LVy2hztTWWBqDirjRKAfmEeKQXS8StDcs96DwFfAG57
BUjW/5hurjR22TG/PlYVIcWs0NChrZvBcF4qNafqDdYBiGF8A4VrYPdWvND8xBpXAe95VSQ47rcy
WxGx03eszLSoGxw6YAkhFpFr6zkZFT7QeuQNWRmvGHKcy0ZxRgYG/c9mRN6NVMsv9+zjuTs3nrGw
Ut1FAHw+83e6MgK0TTNiel2slJnay13uGMGIDBz1Vjr9gB7w5JtN6pUTkCv1HVlLnrb0Y/btg46I
NDFkSg165zBDsvjnlPjGxupwuCf1JiR4OcLZqFQ/P278dx85f+9HgAAt0NwqT1UC+lBPAlhaFjB2
p3H8RnNPZIqyyycLbLFB9Y4JwudZ9DLt7t4sBFFqpI7M05J6H+10DLEu3T19lp1xO1vX0BssRkNq
n2UjuAtVfVEZDTzA/vteKmC1kGIip/jWJN7sCoSNVPqHidHbP69wh6ZSCzQUdvTKLWauHSSsu09W
tvgE8gzT95CZoTKyLhIQe2Rftcj3zSMKlP9PD5Zwzo8vws+wV3W94B3i4GbixtpAwpVAtm+ZnWTq
8w6IxvgZiJ9nHp/popnTLkKlxs3zwg9EPjmmZdDKtljEh+oTWptBMDtqXFPjILwr09ep3nxTr1tv
0wNL2V+yu8E8gTtytsVhqdj4Xt5hLFnk5tR0PTDX6GYneSaUglwQPzIyOKLYBK8bZ9ovZjDjEoJO
VG7UiSFyPDGf0XBfYshUgHAjxK8s8+nP0BTg5ifNqhQgh1mVAyfHvaBkoHtirYP/YyX1k9duKtpe
OkuKk1Ewob9r+GhOF1dutteKRv3fVCFCi03fGt/JnndUWsi+//+2XKHLFDL+uND39HcWNvPyj2bD
uxFINuwu0YLxNUsGEgnkI0FClKVVEouqmrLOAbzVJ3xWS4u1sp1TVJkw7YXhYOL1SmXKVHpNFhlz
BhSWnXc4N55y1w2PoBFwsjDwVDk8DOoylhfFsyqkIwaWwhp71kcA8xUGOTutVZFRwoA2osUPbd6g
vpYZdmwsXSH7kdNsw9qqLm7ly86te9zzHnsitAimBUztohJWoSuBQOtS7AiI7aDBnqMN4k1oeLev
qVRU97pt7SVLzOJ5xRjo2o/Hx2i1qjy+S9YzEjfN3alwG9kR7oSnY4+r4bKCw506vsiy5VgyjaRG
XCZ81ozR7SvYPbCJQTMNpe4vX8bv7lDh30kzql4Tgjypa3FR3my5NqCDgdebHrzMMi4OidNoPZ7y
5rPacnUwLssn49Ngj5eVu9O1+N4HSqbaiDidS6PQJa5mDZ+zdO923rpkvnGg/eDINSTrcrcjey0O
LqBWhVZeFZR696qFXGNBTBi1MenFGRwWbKGrE3eXh71Bdf3FmxyxCq2uIpO88CuW36n+Sksd4rOf
i+G8e5v5a3+jFJMAbcNn8+an4s8Qk16h6yXuGRjTKpZEgbmD7bLFithVzBL6suWr7v9OGdoF1lIk
biHmlcA6yAkpGTltvt7c9gVi8zvUtS0eSktByK/qglDoRaxXOiPSvjNVnQgXfWUQqc9tor82+EyR
s4ga2/4xBigvlVQ6RbNAuFB5AVHJrZx4GSl69CAma/qThbRBI3OmNBAmziZivC3FN7GrYh8w0dQZ
F935XE+bA+19X1tkEvu60/IFd7hny10iqUwe8E8ZQ9m8F8+uTVLaId9QLB3HwkfPKytP6D2Z7i0L
2RxxjBj19OVKZreCxJw9bbxvZJ8dtceLg9FUskQKV8pS8Jv8f8a+pQI329kdllENL3xwYbV2J4Yt
f4a72QFxnpPyBjfcjmlSKvCoGzcuUDNmhWFA54M0ioCwy3UJd/rGNkdbxnq3OwYAfstMokNlCkR6
p6j7gvCGI1Qi1Q/jQs/TjqFzOizY7cITX9hliJM2bgAqJVf0RYsYK4+Jd3ev1zshjXh6XwNKYrhf
a/WvtyNuS7/BdK8kR/vsJhC1UtDZFWlfPTbNHQqNbpIfHv47NXqDMRhKqjczMkHbbmAzcC6x5Ajx
2s306zH3pQazk9n8HRmCMEJ5S2yRoZ5MLwhM/Ovn4Pc0jWwNuL+EIOObAJWHLpgnIi54DL+AMomE
Yz6vqgdDTN5l9Behv3gSiMJ6DtaJizTJeZy2te1ZBsbm73r3ZavXOOv2/kw0FYYEnsM11zc6lqVh
+OGCG/wub7uIrgdiAz1zThbBn7MWttTxCIDd35bU/ItxOZJgMkKo35kf+PoZmGTEeTXYjSRQ8uz1
Y8U2S3aWRqwGiqmY3IJ5LparCOI15qAdxEpVb/F3MgKOyK/y/U0eVhlo6cZ92zjEd2WlpaznnbRV
75qUnL94Nk3l7h5A2IZW9wWWNLzPIAXjsUPUl/8xMSuY9+KrA2L2d4d2NolxDLHMaxy7ISj0jk7F
OD/bpqLQ+eIBxjf6zn/E4g8+Imd45H5humBHHRo/GWbR1K/1/5FK8XOHSUuMqpAKf2qdalSXZiuo
3shx3gI6kbSjfboY4gJZtIuEQctNCBIb/LUiV5ElMIylwdbrgs+fYSAXAAUl2DFa7WYOhcVFFIT8
pdgPQmjMb4NID8hgb2HnuK89Gk3USLsIV0p8RMeP5T7+WP2dj7+cKraaUpBnfi4amFZbZDGttUxx
EDVNehi53dK2BgFQ4EfGfgnWiJNC7BhQ6u/cilHdI+DqlHu9I0nbJnPg26Z4czFEDklwgxz08BJG
YeOB82fhi6lycbyHliOd4mYzm24JCxfX3LvKL2sy9oyCUd/YrJ6hP/R0c3xy88vWfGETcR91hdyw
EjuCxiSgFH6g6fSgE+5OM/Wh4sBAlG7yh8ul8wU1g0ITqs8bQEXyMo4t4EbaiL2NkKFfmy1M5MXJ
zpQZGNqI5GhYCIR6b9+7kLmVIsnihQTKnE08hYQeUmKB3pI9vuQ59oJLmlntg/gXiUIm35r01pvD
nkyWb7kmc7Kk+fiKBNityra2AxZMySZYASKl9QqpNYBDeOcM/JuyUIBnMmwbJ1VZWuG+kICe+sMk
QXGkNMo2ZXjGQQsl+ufBBudJFzJwPsvoaKpMfiXvazBylcFML/HjrIkuYqlmDTCvC1s3DrQAQZ8L
j8bWdknW0R7NUKEymvp0yGjtsYpnXGxY+WLSuBJzKD0jfgRsYafkxK34iDZun5KBBuA1+gnt7Y2o
OBLJqAfI7q4ePRQRHqzjQpi74hpchMPq0bGOAiA+rhHOPEJYORotHGdkDE60P9fyHI28A/fsfl5Z
8Y1PbHY5n5y+/9RoGMcRVEv4CpZpiWidCKCPMkKrevSRhpJ/Gzcgs87iQyW+SAuN/4ly4KE8Z3fs
DjKjqGebZNsOBIiQ9/wTh5GzAt4SGxbARdYNx7L5mDu21etSBeUd465OgJtkualB8PgbFiQAouFd
HJ6OJNOHol4BJn52OzQ5y0dc0zjueMZ9/nTkRSp6Q9z6z4q0gADW3PDA9BNQ0a02glyF/wK5OM4Q
QxzTmnQc/6N/zjjekej1M44TBdRqStte7kDPeqipMa/Od0Z8uVoNvXDQ4W0+NrOTPPiOv+ZKKt+l
uPXtp/cEW5dBZxTAFXLNWxt4x7CRjQb1LnBPSQTMeI/skID6ZWqhhnOj1lP39bBHzQjKToh2QmX5
OjljIdxugcb1IVicxFpYeMc9ZYeGOChzE7HoHMpRZuixe3gJKCI5gO6Kc4hLkSIN6tYnuIleDwE9
YRcRZ1693HVpre/o1vAk+69XtnLNJV9h0XVREDGMTspEGFwOJpUBXqs+ir02xm6auklY5w9aHNGD
shKC4XrWMalnk5I4FZorGmZcb04etMaO/eMvZMutp0fP3g4Q8RlkrdftdskiPFGF6lHMd6B1jAlX
cW4e7VvF7XfrNZFp0SOw0g96rfyi/2PvlAW5AWpjFHAn3RlaepDjCVoeSorbsY1Y7LPbR2uED0tj
3puMXuTZFaCeGRz07/5e4Nmg726/R8ZbwxLJOaSNV9PyGVv44C2x/GyaimFi6m8Y0xiWo+Ikye/l
/YP/m5igi0Ye2RpyjZeG2f6JgFEJ8S2To6xKwRCG7UHO1bnzivibobxyn62X31T6Y8ZYSU8hhxC2
tsiDrG9w677mRY9BNS8r0wRMPptlu68XcjgzF0qHW0fAXCugdEMH0wH37x67JCzXJZ6gt1/ho9eJ
7HwNxz7fg0fdhAn0zbHFDkXG1DY/ODDrmH9OeWbedZ1nCfgsEMzg54dMdLmUQlKYMtYbRTofqjPV
hm+QSluWqGaHVYs/1QiFpRfhIEmtCC91KkPmu8veXWuO+UUhnTVrbzkRTxSbYhtVVO/KuDvd6u2h
k09kYLAFr6bujLx9mtg7FjFqipxbU/4/iJrUEjmqvbMfqI3SFiNwOtul6qCV20qAujTjuSh8ZKrF
obIKddcAPofWDnHHM2OVigmiIstJyXBtYAA1vX0LGitvXLA8Xfn6lUGCU4wSfXSHIYJcVT8YvMQP
djXSaL73Epsk73XcGWgZ6mlpoaCk1OVpHT6Ghr8WJOW7JJcum2azDjhwHc5JeZMp0wt1uwYfkb7e
1pfrp247JfS11cDo3xpT5GVW2TTnlyQITxc3xajtoijfoJcu1L9d3WzgaHHzqt6UG7p3ZYBw74vx
u8mIcSE5OLEqfJha64sMXu6nhIBSpLNEKqDnRRXeP7lrye8xkBhDhtMRHh8aG14GjFJoEEhFokED
eTpBtpNHjaPPyina0U+0xtPMNsvJzk15Dt8olI3lwZ0joBEnv6GlMXWIDuqsaaj2+51+fLpwKKdB
aYH6pTrH/oD5K5d97VH2ulLACmWldwL1BAqfhJu2S6RkAJpG5DvmTyFYEo5KlRgnWq1qBEDLHuq+
zE6eZBt7af5JSjpSflS4SvchOZOGl/gzGEhXT69AwYQyi0SOyzeLvHjeMl5V6UuRAMzvm6l2/HOV
Sa7UkI7shgEb2I5TSVPfhdXz8/L4P+/yiep6LatnqGhjirXtLq138saHbUQSc+B3vQTzARoxiHGs
pSd/hbsHS6JxgqA46nwT30OKw9c0yKXBDJB3g3X/wnFsXlM+gA+GXsj7p3MmHTh0Ec78sX47o7b+
GObVHMo2LStnm1FqVg5xav0cvW1uiBNwhCmSBA9D4ZwGFIZ2qTVScpQafMvdDmCAAWEKA/5tgySG
v4rK/7LqP03EoNgEMbcE2yyff/f46Bqlq8PS2vMcFIqCvknOyDyEVMD/lg53tMbUN2g7vagHBT3Q
GMruXiDnYtMcEtPvb3zwQ4wUO+enzH7a1FxDVbEryA4zI7yZShM+bHsiVFJMNwoTWzMfF+I1YFBN
8mYtZ3ubKX1iiHpmQHBm7aiJjKWo2YobB5ZgZanh32COVm5FdvByb/ewmBTS8MtGaL83AIrcsaG/
AvWTB46FFhqFPM4MuILebZEohMmHyuwo1BZjgR4Jf2faDnUbyxRnVyCiILrXU2Z/KJnwX0DMv0oh
uQMAJzUt60Ta5OPTbYUyZF/RnUUOtQ6CTyzw2kUZzz/fHS6adJdelLln7Waf64wo8NUt+Sz4HV/j
AciBu7oHy3P4h/1evFCued3Lc5Yrjr+qURMnkd9Wan+O5U4h9xaII3b7CMVNJkJYfuewV5zJ1zFO
vSLkhjrqczGUDEB8C8R+VcXJzb0qV0riuA/w1aAr2IOqV3s+5s/GgEH/y/Ake45/zw67my+30MOq
N06pWNs5ei0x+1NP01DVg2HD8cjcHLqFLnR0uVm+pu37x7Xu3rQ1e9P/mWkdzJIge98cs2oV7zP2
D8gsf2y59wWMKW9QSPjPjY+Fn9kI6cXZjnZSrHQ2iVAwlsgWwUF2wgTKbLh8VNAguPaX7SpRpyuB
yY5pOouZ7j7NRdiDbkX3GqpO+zTqDh74iL/OlQv/7BcZV0Bo8grIkKmTNhNJiRgeS6N0kSvKgem/
7MLDMFdDdjAo1E58Xx4hSjJx0DECeRclLRy4piA2m9oUSpaLgbQ9X2C1pUyECgo1BOrfV70skRwu
6uNRNf5M6nZMEtmgmOWBXG7ZE8QXdC5CEdmXKbV4o5ZkhTXi4asBru1PlQgDxXnMsS4ijRnw+zRb
qfhliaFcwOeVASFi/w0xUELpuSkcKbymESb/ujzTWzyVk+pED4A9aR2Pk6rALzLPWb7P8bPiN+18
0uUKo2Aea4AUM5gNfnUDPDlk91hPEmzzFkIWfdombA8dwSoZS07+laxibGcuuwqCIjGDddxOj7AP
neeHS1z7ikCxCw3ut6zHM8BwtHRM/OvBYbyivXIMSRsvVp34o6ldSNs3ljzaqxHJPdXOloxWL2jx
pxNuSvzznbnH9Z2js35oFnFoEdlRM4UzX2Dn26VjPrMVljKKaKqb8rGr2iDW3DkmSfWJtfl7nyuo
Rwri3myLqAW1t2/rE6KXw1JWLNzDR7Y0UwX1ZW3RkgTQPkaiKHEsWDYeaNMJszvi2X6v27/dWrpZ
0gAy4opTZsOunRqNyK7hggD7BSaL2H0kR1A5RaUrbHZ2gOVWZGhBgHNRrqRINpfeF8ZGI7qwIIec
Wk+endywu9Tl3z3pamurft+qYTr4EOmQDbbi6QtHW3jF2ZqaERLbUrHsSnwpSHxtjOunSu4wF75e
ZQ/m+ghIBacYbewxnJe5oeaxuOOu6H7BmDCCu0JMvhCHhQP8/h0qZ6p6+LOgYhupvT9eV6nyn//R
0ZG1QSzdvJ7W3NDfFkM/kx4nh8O30nBjPGCGSKr9EicEQoJmg7ah+faHLqG1bjIBphHLbL64It8C
o6suUjoIteo7nOOI6VrU5vxkvIKMjywEDDHLBxW+3grSco5DxNkxx85r57GFRAL+VOAIJA4ruTXu
ImJfQX3ePqv4jrcFbFwYCWbnJ5lMN0JvV/zJsAyTGgjfUUHsGbF7AvBFUqMhb1iNrAOY6kH39dnG
h+08gGJKKXRz4N/QKd+oK4oULabpHb1war0FQZQKPAMuuqR4JCuyo8Yy+jXjPZiTeDvClpL8MDrP
Hou5r+adWQKxKTqgf1xCz+SctzUlQpHIgVbvx6DHHIMOn+TdaquolMi1muGzlgfN7s9RGFQiX940
J/2UksSTmvXeHqNNp77K0U4/02w8nlPSc3Zn276gortqXPg/zNY20T+0TcDuSRIhnVr6STCI2jyk
53xRKZPx2/B5Ag/d4C02KPYXY9M58QQ9iv/BeKP+y2SwseaMUeCz+f6L1b61of1gfn9kCmMJ0jfR
YT855OfD6mCr5CRhiW6N3vUpiU0Cb3AlDLHleZP1oa47qqd8KniZXEBAE+pEwv7Cq1j0HXL+9bIh
ED5PzMWp7gbOqNvYiJBp/1ElLWAWPp1cF1Vx+/aGh7gVAe1IWvg9Yy1o76r/e2VJnd2/z5xpHTsu
Z5CYTrCFOVexOt1JiRNOAKrkiP7N6sc5WNhADrP+I0ZMQNtEcD9n+5vZRKwL4GDuinSIw1pX1yi+
0e9VvRDKZppn2sst9ZWtyWv4mZBYd1Q8JV6s7+u6diwhs2bx1DO8XxDeul909Ts3axpzGM07aDQL
T/Q3jpj2qWCKvFMeOcwx8uXqtKP0PXS9DIsGlJ61IGL05jCnaaS8fTyvL0fEYMkmrta3KMZbZX1+
ldD+W8UavhMEuBeiPjh4fiBQZ6r/IMb1hfdwfk0Di7B8SREk4Xoh9ejNXu/34SH7dPnnbNMls/sN
2ZKrpQ+f6KUoh6RkXpuAZwdu4BpbY4iPVOM7Xz43O0cF2KBpuva3GBNs/EqZzfxK4xwUcaCwGOZp
jDKVctaewC6USMxch078g4mbtEnwPUBIz+D2n03fxqgS4mGMaTIq1lqn5e+EdA2AS+CJhUN3P2BJ
HTu56gZQyhgbjmeNXlyiaSJLwK3Onhcn86jxcq03yl7GC5og413mNu4/7AjnlrOBY+WgrMFR+E64
XR3l0tt+bQjPptfHO1003a8c8xLtJ6aSpbDREtD5ELBXJmAYbM3ctBZW70VYE5BrgIyYgfV5ZF8R
goeqExxtZqX0xcosYsKYELD3Hznzx8dvSVqR6f5iAHj3eemoiSx9pXqsL89/1L4wCCNTlwiEKSTo
ThLI1LJsa1fOM4cDesmZeWR5eWiOXFYDDcCL5soTZI6t7WB/lMoKDGTt2U3npG+KS/UUsavct0oL
rnLE+z9TdoPHNzK2OvcqKDa6901ZKWlORg3jbxIgM1B7yUYGf3QPvkswmpC0tyd4l7bXO1UhpLfp
JjTLh9AwexzI5cr4zZ5Z7jWhwbfDMD7EnHngnJWVUvXc8t7zgDTW5AvZZEZljTNk9AH/l9Oan45V
4rFcStN8Vm0b/R+yb3xH4dCRNRbaIqcAIEH0a8FGqw53noeiNqhLtRs+NBjoPKuE0j0ckGMPLrhh
on3gjweHAtjDj1igg5Gz2p+eu4Srgas8HiqWfgmg6Vu6Nbfl+yjeMHP8RgxZAfsIsFyy9EHobmIZ
y9hgEAAJTtOZHk/7groOm+wfQEqsn/LLi0a65/PlgNg899wWOpy6hSyzIRKpESk1uEMwmWT88Sa5
uA9A59kG/lUzBIXzmevfve/hNFMs7cj6QvG/6Z4Rvil2zGhxtbAYACnpGJkDauUyj52ogMdqbkAU
Y3aW6Pmdg0/utQQXQRUs2dLTp8IctZwzYIJ7/UD89gSbGSJgmphhLEWWjUmXGOGoGLuIX2kIEnQD
V3Pvq4QndBjcRr4lnqQsIGJyO/cuYQDvpc7PnH1rCkPdml7yLGxmZMGAFv/3YlGdWXxsq9+mcalk
V4dcn333TmNw/ozUmX2+J8vcK1pz4WEEcwEj7cWKH0tNFFVTp+47xynXv9bMvfQObOPdJajKUNGd
4HFgZtZyaBfpOVNhdhvfcQRO3oOXvhG9W9p+p8mhQQCQnAK5V2CplCPda0sgg1Glnh82OMvSLMro
rN2z4dfFh8FxwxuLgLdkn9tvRIxHzTOeJCcpRG/7S1WdPUu8jOCxB4iOR1cIHpbiqeyfZKCbv1O2
+Tyzir0+itQjPgwMMKSZgYSslL99s7t/LopmfAwaoSPri9Ypgq4txQSjqNttEKSq2NOhUzQxX85n
cKUgY/cQYPxht16hFgOO7FoKqnTZmVLIUmZ4R+B4acQ+2XyZvUgw89dGRQYEuuU9P44+fBNuBRfN
jgFSz4qS89P3u4EB0M/3ESSFpIYN/YPkrGH/qJp48qYmf93TKRwBMNBf4oqT0h47ebjeqon5uNFw
q9wpVuzTEiy2iX/niXzjCI39XAlKn0bnPFjHtzA9oEug2TZRw2uDRvkug6xmZNg21WFAjTnZZWWU
gr5vUrHKTIMjzRedGSwY1hB/0QElZibSBRzm6Ctn22d897NeUznNvkpe8FzPDEt7wGZq5iXJjnfe
qy7aCD0f2PvPtehpz4mriNApNL1D4+mTzVdJ5Y78/XkZpX3IQGqg3X3TQCNqPNVl+tcHyCsJ/gg9
gDrCPLO9vUP79JsWrVTECd2YvVGC/mY895f8iTPn1Raj4LyAKeHRObrphObGJc/2CocsLZUiBx1V
RYO16ueqfApNI+eNQgO2UGU+iXJgcMXzrhXWPLfBHUwP/S+bjuzg9r5/8AutKz4akm532YI1nBOb
Xw7VlbZMH4rY5HGdOZL1edUmGwKQy4OcWMCnzFAXE4jtm4k2NmHrgSLGu5Tw1iUgMU10rf0V/vxC
0t47LSRTyeX94SpJlKshgR6ysh8WXU6JqEqBnvfFZs06b0TE7NmWGUI5An7V35unihCUZKyxfkgE
BHWaJ2siKnntdSZXEL0ziTnxgc3UyUKOgGC9twmW+ZXew42dt/T+r1uKEZXGykX/whr5BROxaEn4
ZrgiSKaGTHL8an7sMwpeCRn+KmOlIdDuojrIRaP5dmtKRaoU7/DLNbxttgr4MZBbNaU6M2MZruFg
usWbSqMoxdMbnXeOZ4LYqWaWZwGXWoyrg6l29Wu1OMVQ19o708pDs0QFIj0YAPLTjr7QaogpCA3t
1YoX7vznOZMCS41R556R0q3x/uiOTJ7LVwn0CMzfFk2bcGb38u3JBrS/BwraSgvUkDTYBcJuxy5z
Ii5OYVcGIa18UMhXltN4edcUyaKOwU2Jr1pNcYVqBx4Q+yIGieZXk4O0iqp+DrTN1Uoas5MEWkKU
Ydv3I2Pg+941OHOuORVNARMN63GOeJPVTCrA7CpzQs9BMDs4zQmWXX5FYd5Yt2vy64EJj7hkkIk+
25XcfeKgN4cJea1gmk9suCC5Cs8rSudzq+Pne2NF4ALNrH0E7WAee+KrMq3/GY2rWgB91PCN0oCi
ZwI/PEK2DeZz+ripoKwh7fuvaYk2GTN0lAE6xZjTm6qXqJnbpyrerQc0o0cJ7NcxDP7UpN5EBUiv
zAxx/KUY+xZhYS//k5//Jy5/A5MB2m5CN1/5MZAtlpyEqcmtlAM2AkZYK0ZtDIHwzL8wjTp2hOWU
B68PNVxzJ1e/9dLkJDHMqv28+xmH37noIRFwoqZbtI3dsXm+yGjlBXTMSPpVLdJmXehHIeY2E9aA
UsQffWN86AOrJxVGWJmSHKWx4aTqihqYIwZU44hWp2/YOO3zeQLTpCXIYzvdj9LIqA4HOiDgSQb1
kek6l9UXdeczk73nScF6mCZKOWL4zw+CeYhRE/T2LxgAkQ+mR9oxWBgtsrOgYtoP0t0Te0t+Z5c9
S4Nezn4WvWTHY8AeZZcdVRBVO4GChMPhjincerYbGYgrznvYiF5rZ6Pn5JuUDdfj/gi14/xNjHI4
Yfd9r1iRXnrsBNSCXh2K8AjYDdd6o4F3+OcQwyULk1lkU+02/CSVrFqvapyNR0gK3wuxIFX6Kfl+
jnsLeZIAT4ppWBm/SIDtRm3q+ZhgIilsbEv26Bj/uUB03eQyBja0MR9ifK2tiHnve9tKVpWNywHv
dX3MQV6DgY3GA1ELKRLBPasRCX4gdp6uivpig4CeB12G8R6upHqO9rYlTNb0HapGbo3qoIOAxu3d
yGXCV0jJ/N3pcAAwjgu4Cn5gO2Cj+eEMNk+sLgAuXf/I6+eRyTlwW44ERtWwN23USpP9JghIdWWm
VvzmNcWn8iVCppajUI6LbLfuXEqT95bzHv5GWaOnu9p9MQTPZ/eO6/eWt51Q86sCMDYokEq1Gj6d
aV2b7pF7UYUEzFFt23wXtTuerhFl8lGJNuXQHLCfiL4o0Cx1oWHLHIqoaOf7Iaxt9yRwfjuvwjtf
RzVPrEs/XxO5ie0nhwHDUa9qd3OcypjCsWkcPGkOWIR6qJQQlZ+y3oWnmA6pzusj42m0g5O2TVej
s4ZVwaM1150692eEjyDei1/kbteppa6eMfCxHMZ1DLhmhzoqKFfS3o67qahAxh7aQiPUCGyzwprG
V8sFJ2Kid/cy+ZI/MUy71TywZrogItpMoHnhk1/LODWkshISAixFSLH1wD8dDMR+IVHHi8N7c57f
VwpkY4Emn44uIZgJpT/5vVLgpOM7JrZRu2+HQktqUjLzM5qYxmDlwl+CR85lL2y79anlmJbfMC7f
HgHcVzikwjbTNzAL3iyDYnlIUD0e34DAHEhW1Dk2C6GguDB5TQ8+C/8gvkVMz5kgm1Zo6CvBmNYP
8mm4xb67YLGU3Z4AF8bmLvNB/XrvA4ZLh92AKToIsoO0eCf/2GTwtlqxCWvnBL0CdxtyMAmR7Gt+
5ZGe93ntR6rditbOVLnlB1SkicxuABidvEnYXdJK+MHGsNqXYY5QZpR6/hzK/czHSvfxAI9BXyKo
zXumlskDqqxmgjXD8KKzCksCTwdGmY0gZu4j70gOOhi0kKqr0kLb+vIY1JK0+m/s5l3GmcFIJfgu
VVeHbjhaS9XHoqVUuNgtjjUvTf8h5Q/zzjDIZV661zPkTkKDberXAXajwx+ZXSVcw8j+pw/7uj7n
IQ/NtBxWOnj7x0/owgPZ2WeJSpf3H+1CXhS5VSDgEMfQJOgj6nspNx7gQK63TwXFLxmbJ4kp34tC
5yOWYNwxJPejBeITpjS43/9SohBBL21oXqpXSP6cmQ4dyQytyZClG9UG0sJecax6cb3P3Za55wrn
r6KCCuhhD0caYv2YmIQPS4Yx4izwyxJ/dCJptEYhvB9Jk4ACEnAii9oJgqEORG732M0qxs+6a60F
ulYO8qwMoBKkn/ktp+gF4k5Qm51DUjyidu0iR8oKOjxT0W6QXtMZESYBBxBU6Fk0cTCEf2IXiySD
5tg5iYZ3xX2zHZGxvxKkT0DmBHnuOZ8Lr8nZGOq8TCgApfmxeb3FnkhN0whAkAmxvkvGigTzoqWB
Bn9Fvg0In62Q1HtXml0hvdUKkn06fS5Ndhrkz9UIfVUsN56sM2On0aCXYcOl1uviAtfCfAVsp7rb
ySgM5jKhR/e0+dUOmPedszhfuGxxgoW8bge6Mz1Y7ATN4dqHL2LOXGfWUITCPJi5rNjWpnQzVv0j
5vpaOYMYnWXv3hCRQxzk2FikqQC11PLDZpqvtLcnjGphKgks0g5kcyfThKp1JrPtp2A+8ym8h5bn
QdHE/tKXoskV72mTmeUViokjzhfgrmH0YpRDam9C2htkOuJC7Bjd74t38OR7xs4mewvpLBKu51tE
ruEOdbTH+negzGfhW9LTXeauLqZdTpP4cp1c3n+fna7+X3aScqoKwpDtIb2OGKw6wnIK4fXsgzg4
wG4tzVDyUgNcvnnTktbdYUUEGVrfH5k+wQJsfYdKTTtsQc1EBM3BC5Ql3p/Q/mfa3UVtCZdSC7BG
4lM6e9i5SQ+GfKDDXk1yfT3vI+48H0gKGQMCa56JVXsz/VS36G8/GJfrIpXwcvwas75V9iz+DGSw
7tTC1pWKm4TXt8rX4CYAkWgp6KVlKS0c60T405Ah0Q+XcJRLlI9fLVxB2LSk5lwDqWZyv1T+Zmny
96f7ZpC3fyYAy1XBnEucF5PchyhLYrBEvIBRHukgJhWN7OZDLsZF2pPNC1KMrZnjvrZrx/vSQVGm
5B7KcVfENTKMw0YOl8ECHJAlZihMMZ1hfDhhosAmEwWAkTZUrOraJjDR8DW5NRarikRMQcIM8zlm
h5YI0Ulwn4nYDvYRhkKWb20o0BG7U4xYXlf+wI94njQ9tgolBv/IFPWinMMuqrzFNUXZk31xPXfR
8oXU4QLfURpIZ81sMQtm0LoLJQvZo48rdwD0bDm+pVkcGRcu2fyJmK4Z1Qey/6sdZds9N1jS3tHM
aqHG9czpvpqVO6GqX8E5uvJK07yM4+oD6/06womL6ooyaeMz9P+8nPdnUObNG52+YghC1VmPGgcR
COMvQikwyf4e6NJlX0VFQBh7XWAjEKV7ZPdm1UJEAXBFa0t/2qNaa47P/QyMf44qbgN4+OQAH6iO
467nVN6ga25eDblY65aCa+SL9364ZxhTAO0RmNEQ9fn1oTiD6S2qmCN0MgzDHL+00ZXdVERhJS88
sZlyUPCZrrWSqb7eCBVlhXLdMXcRbF8z2UnZjvOfiCdOYrECD0xZPw3Ad1dDsxS4N0mfNr01CroM
IA/oaXvEM1Bx4y2XxA5YxyHcTFsr+JjTIMqYMiFuxZu/Bl0J6i0Uw3/pDSBlf7lDqmr0BjVYHyf3
MS5e5y2zAUwnbjXfgpmhKu9Ajswvespr6ARSfw6J4RNGhQTE9+S/NrYyCOI1f+Z8eKj6cas3/plz
dAQ7VJu2FA/jj/9eHFtWw1V+ukM482z7DDWCYon+3COCPhElBkYQfyl8WT31+QAL81tKHWQ/YMNx
Ps7houfvUvP2r+Q7p6/7J2D5ABfIht4AB+4c+hMPn57g7iCke/vVJ6SOe1CwYPL6TSlqctzB9yXU
MgtSti3VUQ43t82K8iyn6IKtIB3m03pZyKBB+XrVRsWe+8J5C8qQYQcydE7LIMmAlNosvUlbEijn
vnlvI2PBEG+tDUlqKE5xwq2OwS1ilp8rKhKeco34RISc+kK63PFDIvCOWU3cFnEAGEBBFsr8kLqd
prWjFzElAf1jsgaeQSPnYatSx91jTRhSQwNXvebtnZMKnMCoPMx0ARrSNxrUSYuVYo/rXeilRlaH
iWhZyerDXpn5wEQF/ugmE7pKQAJe83BtVK7DrCL3sGY7oGwsp/Vc/66tFhMrfgBRGiLKXqeAbx4a
dqYJqqjYPQb5QxaB9SnEZDNfDaZBKbuxZJOn0VWaq1wNvoY6Nh9KO0qJPJ0jXXNmgzxT9g8sMU4k
YFH/08TCFGez28vxL1nl0wLN+FqHDibKKma/xrgFNVsDXu093KvM6JI3o9GysgWkYmzxgp8jM1yp
TaJMr0rGU0QwPGdTD8AkcQbdRDvqwZMSn/DF5k3+md6Kb2iIpVl4RK/lxvdMeTfGlt3VpdOvXpYm
Z3TCaB6HwcI9jukApi7jDF1exjpYXI/ov9oxK05TAOF3zOlMq+ZB5mv9f0LGiNdACAcBIy1Su22V
5qZgXQCyU9Wo8+2Te512/2B0Kbyos8E+JZmwkPJ3cVr0ux8lJVQ+HjdHTNP/yxL5hFmjZAIBBpjZ
r1yjh7p1xZnclpZl5NGDRT9H1SLi24QY/YxM24iJp3h/laSwK24mbYYHdW4dgmr2ZZqp+s/G0eAa
Kljz3w4ZQHAGnpNVshWn0t9X+oQz96VqMP+b5ISdt3Yyi0C3ypYz960GsFVVri9qtX16Z7PhpsU2
tycp7otPjhj+13fi1rcVgnFtUDqeT/XZnOqrtN21yCEDFk637jXHAn5Yw46OlKv+xsV10UUyDdBM
2DpemsS+ZahfgL+prUFx70Z6dQiXHVOeKXPj5M3wFpYGJ6Hn3EPiJcAVa9MliI4gEsKcwjbdfjm7
N7ezxTLW5fSMsuMzLWBgzMDWNwjaDRk4POwBNcKoVutpQy+341jXSDmaqnDbNt2F6gmo/tS2TbRy
v49Z/MPlG0WznUdIygAJXyV9F0dwQbIDocWMAfwSc4uE3WFPGsDqfaxp/GmFX8kzKS395zqfze+g
Te4IJwzVjPjkSXoRlWT0YWXEXUZj+3lCG65JC8seDUZFlDwu2/6SumvOdhUFFhWfCrTcc3wlITY/
vKRv4NZ2HwJaQdwN8R6n79/SMjdBxnGwaBYhBiKXH1PUxK6vnifdXoZIzdam2NRFXu81WlxNIrJJ
YBfVoKF3ftsXV2vnxmEgJKNXcB126mrmIy8uBBWGaI8VhjWNBrQI/BMsaH8MT0tg6Rf1rBB9zlSz
jiwMRG06M96Xe7MUPLfUMPrqfgXw9o2zKpLIojYuZMYoNxiNl2/RfNjuNBItWfdZVDkEzIEeZZvp
YNuGLPtAQzSBe6SrFnf8AaheIfxCPPDjm1nt67ClJBaEFya6aa2FQKUiTArpJ6aUd5uv4nh8lQRc
oGwJXqF0tNUbekaM7l9Vz239OyqUzX+GdgB37xs+VsHmrl0SnI+xAe7ye5WHeBwAUasuy0f6ndpn
bDU4deBT8/18W47l+SlKf6WbIdPYmD/LzMi8d/TVelD27omhXLXM/botrA509rfH9W8/BOs4gKxS
9wjR5+HAm/phZ/MK7N5nxIu9mSgb00ZbGT7brd/UzE8iHIY+0w7PnX/UzPw7BIYwYHENIl8+Chiz
/xi5jLIWfqtbMthpIsbt3Iq8KIrkB5BVEt2a1PCUqmt16GfChbUHWFLsqqAMoyBPGcN2/uQfA27y
iVByWKp7mb3EElHhMH2U/JPFEcC0jzh11piRACCzUhbRmEXnhAnojCuxyP30f7SjyJ7Gfi80fs5S
x6xSN6dat/mQNpBzlkfaiyBARgJK6ASwTlw49zRQN4yWsZNPIxL/aIpmTbzx+phbgwdRZEEfjifU
cZsZN3Qn0aXfc77Xb4VICh5lvnGOXBC+jRAoKuCJsboIy3XFCcCQO2OAbRIa8pHYojHSK9z2DCua
V3/TJc5It4kRbkVvJmjSo/TUPkWJA48szKwCxgXmkgj5OFBD5X4IdDbB5tSm/UckbCdFCi4ruja+
w4giV8uwCLCdO/rg20+FxgJCOyGGMO9OoSPI9UCXbPXWdE2mhwNZs7rVimC7jOamRTcu2Qwj8Lut
d4ZspUZujgIrYHXWX+hiWaZkByZ6gRZkRACRanjhz/bmHvR3jqUMgkV+4KYpGel9f2kcPkrVdwhd
MF39c6/RTA4/Q3hKJTwlMxpibD9l/C6zAh6K1aiaDPMqorRdOSRlYc02nRPUd39xFJ9jlPtLcnwH
m0+pHKlSk5W8cb+7fy8Ypv1mv4Y5TQEAbmiT3ud8nRFDmKBOq1D0ChVAh8Xw0FgepX+J0wyKX+O2
0Zk3nBHJCwtn+OPibL6zpd05Odl36H/BdRPDgzn/W8u0Gi9olP8JoiwAGo6j8V0OgDYMbogyyQex
KXEMPJS4s3AdgllE1N73TciquzfHHGgre7VlTOzPo2zGMydQvIAczpXOC9zE2yDLxYL/64zo4DJz
rYFsMEpDXCL8q5qkaH0CKH7FjPvWTNCLT0LqM8CvNB0BX9JBeOxeL8nWUABIZJNMcsIdyBNssbJr
aDd3fKbIdrsWgVTqjkQCnq4xlRG7UC6HL8HMzafihMHxHe7rfWYicqycKveHg54HJoQrrFQ0rcuC
nMQvKmcaBns2K2BsCFrpWGNWc75aUO3/XAQGR/8xLZGdOPUDh7mLO81tPB+lSsk2uMftSg3WsxJ+
sczOFtd7fZ0oBwINlb07DOMkgxqDkhKZrcsUR7j0VGp/fm6DJP49cT/n+S9B2UTUDqK6CCWgJhX3
FZlvu6d+rLcZkVBDSQLIFQah8bQ8NilvnL/HfLF+91oeMwl1VV4CbLDMROItreWXCJKuW3vX9nTt
pOM5ruyDGIEQUbTeTt7uCH9p7JM6+EWQ+GUN5vg4yVzqI89HYtiEV8HfABP9kJpxrrt1U4aoQeXA
cRSuKzw2kVtFrIqDljcwXqBPAoHtMcV7jVVopZkVOYAP8nLUGbi6ImZwgwqLpCYu1AXGh2VbmZse
PJDraJ+bjUSHr3GMede5IANo23WqgOHEU1iuKlEFECgT0HmIaSUBjUhmxMV5OoOy7uHA5EdXLZFC
tsZv1d/7SrFE1Yu4T9VZ0QJTDJ2DkHC5SOvcXeID+CLBXX9L4uChYm2iZh7QcamP8wS2Nb9/kZ+e
29FcYDC4kY7sFoSZzSVkhQXAgo0JC2rBrD3v4SWIRNwCCPPx4H7NFUgpwjZw2Y8kvqywJ4aobpCN
P8apX9FySFTrUfvtzBrP5ULe9hn+NLO7jxDqK37VAgtRuUj/Ts0/N2goTK3rzfOwc0BVib6La7vF
UJVD9e2mwdMeNwNL5Tr9wEubO3ZQ29HaQ5XEOyuLksGR3zGYZBsfCKuuiGDb2Gc/PS4puInavRAC
ythFpWRhul8SPBeqWnsoa5yuNMjUYXENuxgqYFEokr53GjKoO+LmYio4IPo3SoUm+Ppo9VFmwYOt
hbVD56gBgYC3EE89GoXJBPYAqZYbLLM3vHrta8DXCWkuni1RNJqVaIX/GAU2uV4ob6V8oXoVJViA
ep5uhuE1zEn435lqSze3D4HKQzaw0x30EhXjm9zc3Cp86u91oguuDxvaanuWmpBguGe/+Wqddo0h
UCGFODsG6r4+MXcKSSQbUEHCMt9EOYEWqzYh4BrMFn+tJlvEO8kEXc1Kq4QJv/COP8pTfeYEHjAf
exbjT57CBCvItDUlZbC7gOm35UVuYRPU8+0X5Srb5Opn694npszmzeNzDu0QdgWUS0UY3rdM+MrZ
2d4Muv63PLVpOCd2FO8ihpFFcjav9Fh/dnWjYLALfmGVo3c1FtZvSA+6jJkfHIZVLhotDkw7HvHi
JtnL3YkAt+7h2rNGxaa6UEElnyX4rwPnqSpFLnjgTMyh88mDh1rdyrAlNOtRCHavuDuBGBG6K57S
E0DaOEhTKlxsPmKmCZqOBLvN2T7QeWuYJRQX7CIVx17n00GmGFyo3dCCfY3V/aFDf7yxE+kBAzUE
ZWdOIK2/yGTpJ+VrTRV6BaFo5A0NLrXDLo4In26ZmDXNqDe4skci7KGTDBwnthe1XCe6ctjGC0z1
98Aw7z1qJ/XqLSJuTbmklW5dtxySFHKNI9zEqCi9KA/9kD73t6MxtWQjD/eaIS9holSYqAHgsZLm
BMXIMESEW/drwvXACLxADj0H6cFNhi2RD7152VuP58U6odJif8/eOLsgKIue/z4jG4BGPylQTdk+
TA1ioBuzHUq9U8Ps9s9uN4EBHpgBEgDGEqwRX3cK8PNkbG4ALo5S1gzmKliNC6IZiw8NyuIFvC8d
RIrm+bhMBcOKZeLDhfmADG0YlOd4dLC0f6z538WZUePps4Hactj1vgrU7GWS1dS4OLudtjrR6QoL
Ro++8YeSIi+GKrajFJkEgIANwGQ94/8nnpSW49PevKn568WH5ltMz65Y7o4hWxxUxWhbNEg8f+E8
6mKQePMrdDii6RUFWyd9bXTNHk/SQcyn2XesHpouRqY8lZrnPuScEdncTobBTc0vxokjKkFRmtKg
OhXxaZBzq4DhmDAijDm54JsKoPZMpKYGL+LKh+VTHumwjjqJe45f3MYmlGQJdks/ehXA6oClsZzg
HDzNQzW/BFAyePP/9nx4b8Cmc//pHi9nPOiwxWOihe8bA1u7itQOX9WgE3PnkbezuHf+RY9U3YKD
phZssjpaK7ij7PNqhQHmrnyBuFJlE1gsgVjia6DK4GygheeiKcZG4xNbmoV+F52Ooy9L2RoPstMY
B1QbpTvwfmjphCGJb2IJ4+UOAajjVHq92Bp6tMQllglSqMhUVjH/jOQ1vQnj3QQAdV+a6cKm8kH+
Th5cMgw/McFE0UBcmrMbpsj8gdVhuDGU0ZREFy5V51zi1FJuRe87q9vljvQSnxRmqcMtupUXpb9q
P3CfjIFUDQ9eM0dI5MO/T5hs8IVsy5BQ/RL4YMAdlRiYDIUZyLkSB/88lc/xplf3CPDb+Hp3PUzV
KgzJ4lSeHLJFRqPxaUSn1FKdsUz+dVKmOWGbntYwx0RXB7aQJBDmH1QjFw9fBtJVOjmGdxOcUZEW
K76tAwHol4Aeq/LLWxksxe643l6hkj8edNThiIoMEegyHmiMOMDcN/I3as1U+ZZgjP1da7QZXxIG
/TXPtkhC0Kk6LNkLdjjsotmX8niuYty3eqn7bldR9lt1FerMFyHTRFiGjfy+K0t13UAY1QfZ5WKY
RRsf/g5VFvyhcCn1bbn4vIy38OKScgnhvFxB/nceUwlQjLmrbSZXjSObe4DZPnHlYiiupL3Ad+y5
tjCL4PG+PURrIEKOkmXKwk89nLIvvFKtSG5IdOPy0Gu85DJ7OHQuR02ivZ7iaxL+lRVWhEjsR2xD
+IITxLZk4pBe07dq50KEPsli5ff5qQocOZ8jabHAHBui9kSwMRd5Giht2xBtX/DW3SWan7DJ0AhM
pfh+GErmFhfO1mf6yx6LTrxJwb1JsHa720JAf0wUezofxUCwLOakMaG19SM5DYl0ZS0WlRy3xpqk
RKBm4HCvXxILqgWQKLaT5f57A1aFqkwJTcs80S1ax9r+FWw194ZUVGHsDN1ypBm4JxxSexi+jJwr
+/hsOjT7Hi6Hmd1hfBYmXpHylIcr9icBUIBOA698oNE7qhX9nCaDxzIb8rSPmE5lPzJ6dW8JnEIT
zm+Rp3Px2bF80oY2yCzy/UvsKHOCQQqj/drIZajbeJn+oFPzt0KADeKP+RPnb2dL6zFvy5Qga0ws
8HzmUvi6tLkBxblXsuUDWOpTyqJ1rfhB1DujjA/5RCTMksARx74rc6hNprcdoEUkqJb5BOw1urz+
ZUraAkq9lggMiYz6PAPeCP/okD/9DmZewJn1iI1/FyXB+8EWe9ql0YYlxxUbFEoFO0i0/nrttTZM
WDIgrpKHSFKWavp/yrAisSiim09r5+wMRj/YJ1+fDkim1t5iBJN/BCsbjjoE9GCHcGPOPcAhqzIW
J/QlIBMxaQ7l3VWhVDCopz+oNRf1Y/cnqz4nJRvdmBB2a/4ih95xYGaEn/E4kEqBvLlU7dUWhzrr
flEQTCnqvQvJdBWX9lfI6woHwaanAzMiPsYtimfdlu33jGdrez1LUvzAxmuBqMJWSAQygmS+EiEK
BStg1THTBwCaRDNo/Ruo/kknDX/gmvB11OeqRRwhgxehrl2RBFB9V9hnQ+4DQnvjX+uOAsQA75N1
96i6EkJP5s3aK7aa3oxsBrOmGuNFXvwFcX/UPZz+nmjxE4pFyVuwviJ34XrBIfZKgYSSWQj0sBp3
bzNKCMvB+lhPzzX7papAJ8hb451XaUzHYmSMKlx7/aRparD177XLA2M/RWoXZqA5CAEQTmEW/5ZQ
qqTSdBCR1800fdDBW6bjBfHsNMBA7HYakwM3rTsmlXUwJMR7HWvUr5DnlQYjRjYURCL29v0ClL4r
/QGcTEXHU7HaviNEm8In7kyAsAV3KYt4upoysciTds3zyVW+o6EcWEpclc8BQGmG0NwkB5eCoHf0
BRg1hOY/mI8Suo7Q8YHh+dRFVTQ9/knAaeqA6D5zS30F8MrqqvzGLy701pW1Kn9Z4BVd5lsIeIAD
2NMWRua2WugNAvahDevb8sbtjg/mPG3e35G4bEuT5s+u8Z9GcPmOqYdKsfPUJVv2aqERHdjCFxIZ
KyplDOzG94PCQKBK3fwWRqIfkexT+AdXOIML686EWOM9G/+AVOJ2D+ly5VR+XJKMQrY9L4PipSUL
xGdCpDTcOLQ0vEQu03PuiLjgsS80KowmVLFcQc/OpRFNoBZQVWMUOp+ekkVs+IptOuA7tu+3YiEv
mpHRMyAgGWyJhgMtZmf0mRWQ8WOsX++7mre3nsuCbF2JtO5yDLtEaCWGgqhzbgR7+BFa0yL03z5P
ce06QTKQWIhQd3L6Jw1BpQ3zYXIEhBIB20VE9GJQU8nojuL89TXIbfPDMzsnWtw0ZFx0NHRGF2Dj
MNCRLXUj56MvEWvtIzq77tvJRbBTgcbBVoUIVIEiL5cFCFpQV5zjRAluk2bhbHIQ0BS4HzVG1orf
5OcHJ/eU950apJlgVNw66dcJGspYyAGgXOEtIxmv345m216tfldDixz7pdFjYA3vy7fBIcKFFhDr
niI9HTqI2CgK1HK3E143urk43NqynMw3G1aG1omSJ4M18Kb/0YyqLonMHhVnGhlskkocMcIGTZSm
DCilykv7SdXAjxbYlTRrsyUUCeIZ2jA0y9a7Jy8HfrtBPNCcWeGo51sWoRb5TGDmvXxYsqVH2OKM
j0oZotayo/UpYq1gyB1eiCKn8XbsFHOQrrOXvDZJnEU5BvucUcbAyISSo3WK5mF+x6mrRvQ6J1yN
upMM4vAUAXbjIL7Tv8Zm1C1BpBdlxAaCRw+JfKBe6tI7dY5OJkrOfn1Vgvmh4k5y+O48lEbUTyZW
KN5NU3EcZUpa6RjTM7Bb4DmReEIcgjuUtHvnQ57y2DLmoYoh6J1vRZ5n6Kyw6Piz3mKz5VdPkfgv
eQnEq0UDqULTQpi74SeOlAx944mj3VEWjwSbabD2LJJYwNVThMBlinqHbmFGsQ8jwE3HEhBm/wL6
4q5i6yiWWdPQ2MfqjowGw6dFvgrhfdITKwZ3TJjHj4LmjUzPMpJQgYhy0tbNMW9IrU5Y3qUoZEDC
MUD2q+KGxKcmQUHjh6q0UrrjQDaDO8O6GtOSuQUWkySrMHM4k657ipwP5C5l/yvhwzgr7nTOi3Qf
Hnb7KJBncaqP0Nu8ED7lSRK26O4ubXVL0NkG6ZSSNUxZTb67+knh52wVbq/eqcasQ8BYRdFN4trc
pSWqNOyIgBiSw3yWdUaXG+TpvHtW5FwteNNcJ9N4rsQ15Di9OxY6QHx4wLriBs/aACzNG/YMfknF
JFan7vtg1XDyFwEnju5G29ttL5wdjDMkeBzPO1RzRx2svt0bdzF3d+JCca7/KmBxZlXPMqSqRaUW
N4FVQwdhz2j0xRfqlMbIfI3TIBnc3yOhWHGMPgApowcQIJZESomWNtiEAYbDnvYwwsdBnwwuCIUo
27nlGJ1ojJnNwwcKM43w/PjAl7dUb3esNp09ASV1zZyNN3g7YvYpFb1k/k85Stz1kJzbRMeqBPIT
vUUhU6bW53xgQ2MGdx/s5LvaV+0pIPcCH+/B4TEBS8msl6NAutDI388avA3IKFYCOTZlXlrLrTY9
NHpBg2vwKq1prZlGHSVjng2IBkzyhU3qtbMtJGMtkcP8Ps9xZGpL5RhegEOs4ADZCJwXdauIyjIc
zw+SDgLuj+CZEXcLmFHeQfSPSgxIqw3zqlqUq2WbhzZqLc0nHCHRkgfzS+zdjtY4xgYjK/kflnPW
flj5HTivwxTkNJEWO717WtDPDPrOQc1F1RgAlRQWaBHNZvgQJk7nGm8ph7zI8NIAlcJqTKEfYo2l
cvpCjw+evmLQcYPJGcmQAlfCPaEaKbcFsK4D6BR/OICNrLhy6VBB32ZoKoGxoC5WGAjty4RZM89o
aeT43C1CBSmQIdVnt5K5eu9yNlf7Cqh28UKN7RsopD7EI7lI11xms56KnUV/FkPiiQ0a0s+V4vLK
JzGieJWJOKGPGkVtIfZedO2X9B74AW79y/gmM/SXPRO9jU0+5kpbYNYAegxUItrInSlfgRdanQWU
TO+zOb8cKTufXNQo5ZgBjZ+e4NHPYbMPH7qGzNRvJEfaaikSE6gcULVwnhgIQkaPY2bGEH5Shs5/
FVzivPzs5f7GQ4l0vF4L34RL3RAHeqlLTvKvCTkBYYUojh5xwcf8aflbbFkKs+Z76pFwGd8oJKSL
6A5ByCEAHeztu7GH4QmagxmsNEp2z++ZGZ3ylUp8w/t1hQvE4jXyiX5DJqVS8JCZolXs8Q8pZNi6
+5yb6bESExMvI87RN/rvqjWMEqGkqgHseXY646rGMza0M6zJkmuML0naOzBl+Vd/0VPgc5EMgw4H
cCLN1RlhPubUHqdYD+2zf8BHg7bQ1yrLOOwI30YMcHra2lnvOTnknL8VOPWXEjJnQLGAEGDBLVbn
IX5WKvQc0GhiP9eNnKFcY4i32uM/A3ERZ+XiW2IX1m1MGRJvP3Hevj4whSxlPdFpkPkWbN2yAqoa
W1CpLoQicFoRd68r3TTb7P5mVzPHA88kp+mVPgpDhw2YOKBQxKzwzMPoSS+MiMqWO4k63g5r5wRg
OChI1uB/vSHLfBVkEwMTo7uwBA+YQWbwpBPrG2rI7dupo8vvZaq8OrTrJtBD3/K8yhhwvOmRKsj0
5kNicba5mZTDXf9wz0JjsORQ+8wXAplYcBUrHqnarRmbxhz3KHJlfD3eANAm5cpV02OGMadAvIJ6
DjhQlQVrkjjpcBK3EG+so12htCjJeYdXnP0QGHx664ysVnHZAm8totVuQnhEA9iZK3l+3vcYpvAu
4bolQEB8VVgxVEh5AiSSKZ46nMncPHX5GZwaElhT/UGlQFE2eAMBMFOjY78W/wMkTy8t+7GBEBIw
4dIbsb+YAm8DTQcd573ud11BgEKfAcTsfayT4AOs34P3w8yWpjpnWGpgAn6b/15CKVZVHD25YD1A
zITkmAr9qwUXxQ6J7ku/WUII7ql+S6ydQSTJ1PY/dKrJQXAESyQN+rSzS3Knz8popJntT/ktzsCR
6L9FIKbK+O6Lu+4zhHlfejfJ2EKICsyGVCN8UQb5oeVWPSHlTx54Sd65LkIyIO3aMwtrAcnI0G7q
pvW3Nb/VGye4fw15SIs3fjLSpYohM2avpSTahsqKyKDlhRo45QKg5JMUeEdBxPMCQI31ElPLHOTm
MS/MU09mP05XmyiI8/lCeNEFJd4E/7ZETLKgBRN1mJFy91wL3/qaEZDOUlg7d93wWmnW/Q/8fkZz
mUuMB80Zq65JdWw0UKf/HJs78sw6QYDd2zckNRyRo20KVDuNoKp7rAdSyrU+fkhgLGHjSt28iHbV
wrD5Q6BSnesdVasOWeF6Aj+WXjWNk//WG2PVXjP29ZMd6vfND/BCWnK6i0ELFeYAnhE+og3imXrk
ONL11Lkzi8YLjaB9NowjmXqkbE2JnBMc8vQy+YpFPDv4RTWcvKJttWPW0X3W1Dt+Y3GwOEFKsrqw
z81jAkaq8WDntCO22JjZ7Vq16w4kU8vscouCy95hk6V7xnCLGsfbrYlMWfQ/MeLlIbu9mpzNIRu2
cbeq4q/gVgTZFC8OT2164FH4BDq+dNJL8198dqqW862snxGNnJcSFi0LmEX9hBXswaNfwqfnyZvq
APXfqDz6WJOWU22FNU6RU8HkCTx4+d1/xkPRp+sHDaFga4YZPYVpuCYf1/lXBVUj0tArDsXIL+MS
bj+xEe+6kwav8GkTTCfR9OD4BOcXj6U4n24hBUTaYhyCsAL0bC/gfZooT7gcW9tTs5opcZwjuV80
FBlY2hpw2uiWQetgDFAet9zjGCS/5FOJYWTbwMbWb8LCkFuxHHrxnHSSkG7mkwTMQpaw7tjyhm45
S40coquK8HQekIlWAHq4WpQQQ7qIFORN0vWiPBI069yx4eK6aObt6IA7iK/KXLwk9bteSB65o77S
+maUqzS5YL83f7FGtGwiG5mG7c5Y7YSVSYxstJ3KM3ZMqp78rZHX1qIN38Hx+M13uDAYt9zDJeGY
OftbjmlWo8pbYTrb6DGb6bYeJ5OTlKEY+ErgXtJ/HhMkT/+owBzeesNnJaLmW+2whtDWJ5P+qGSj
fP9AIqooPFiZ9QD3wHWZSKUpfAM2tkLmrTgxtD03Vq059fWl21radSV+HWeBZmm4rPgIYeART1xd
OrGWLfORKXQzKqMeo4NLb7udUR92UVvWBA/gA5HVU6pZVkeuDtyXt4bUSi5xNaxT2Nm57jiXLnyd
avO//bAOm0a0Fg5ewljw5bAYFJ4bZIg2z8hNUjA+GxXxzU38lRCCmgc1y+UY2VjssN6/1ldqXYdt
mbda8BGHq2NFxxrZlzYw6oD7CPsiYWXBwuN5Hhea2fnV3mR0SiHcZt/OoMmcBZv0PI0dTDp8FuHQ
95w8mYhAlYjPWu1zJ1RUEW0NWzYHdukKysHlkLJY2xo8WJLOyZ+7/CDoHtLsmw0wgJzV22jvXOhk
ooWwa2GCzVCtYvvYIIG9zmtSTk9xJ/loGQRZ90bYnpomnT5nNgS+8iKqUjKTWfdUjR3cgLTVjnmZ
8ctXsB7xZxjrEuSjP5KG5xs2+PECAJI5dYhZNXwLSiOEJ+N2Pm+tlJg+WtVirNdHp3n9BxuqlW9J
TTYiY3t8LUZ5V6Td4TC+We9cE3psQrhriHLuXn9h1dmVSdaAYKBuROcALngefevlG2mwcGJQVoz+
M7aGsru9LZ5LURzsogwvNgC2H4gM6sjKCeS/KhJHiSuiPeZK90QnJc+vG87cUBtCaXATczIJO1FN
yOsmeHGrJZs/d2VPSHF+Ly+YUwXeOtNui4L4t/Gb2miQylYO88Flk6jp+OWnCtqh/aFQS/10uF48
JlnLgrC6B6Uk9inUVRJmg+l/eyXjyKoYEtkOjzFB130+VgWcOyzN+OUUuKPYfR/CEznPQP2YXWd3
sQJ8MikDqFaEU6/kH1SYV9jRZnQJkhvdmCB5zZe/bCK0vDZaKWgSrXIMQkC4oyUtTEAeqAWcE6jG
EEP1PJ2wXkbXxIl/wOKQxmip8dzfKkry7naN/jy7t7QzMCy6DabmoKLU4zKstD/zkS4AFECndRI0
rKWvh04sKOsSsC1mVoNADbGAFNH8hrdpP4DXU0W1jyX0JNFfqcYASscyq40kTEVRjf6snNl77MPE
35ZgDi0HVV95kV52YWNijLamUrhK9Ob63Ifr4Rd7cOJgyREbNoeUAVlL+zcypS7zDNPpHkjteSR0
WElDwFT/pi+zxqlG/g6nvSibkTog74jUDKxpAmqXBS9ZMGjR99mQxdw3J+4KUT2Vw2NYw/IM6Vfr
mF8WWsXsUtNzfaWg5gXXKW6fNJtQdsqrqCnemrbV1J0STVNsabAVAW05kdnNFeRZ816QT9P3Jews
7Wp7SInF353kRvYP2eIWxd2Nc+QMxjyjiCoEayJLQWSYv2sQ3Gi9S73lmD2u2sCBW4/AybDuINkj
ibiVBuOuXPP3IdIe7niDsTsawYwD0GagIJjiqiCO/Bumv8N+UOhNw2NoloxgQRbsrwmldXG/37Jp
R0uF4k8/ui8fCRXJYkSJKaWntSopgiU7EVErXazRzIVr0QOTUdYofGmgMiPfuaV9w/q0EgdFo4fE
TQXKq91ous8wP0wJIUdK5LTHd4pb7J+Wekn5uDAzUZgdQaa4UeQ3C2guKDMOUdNHxNOXMfSyn8pl
j3w89ZW/DCoR9Yy8xXKdV9HEERpRObrbV/PMQbRpskC600RN3TWeQm2pgMUC/B31XAGD0VSKhdaO
CpgBnQFeMt2owJhwOF/oaDZ0sAbIsufg7U4SUp5w7nomGkM2NAHaDfs2yOu/wCWhVtSdqabzx4LA
/rtg98zq7pMtmAb9bGOo5sZCh3rNduiEN78wFXBD3vMgieAz2dU/Gp7h7XGnsaUjSHOC3zX0IUOv
8QgEjfClOdm2v/zmzBJy2MIvXCiplP0KAmHjS/77al92Ngw0qYDNv+VjQX0yj0Y6+8Dx57wQ3gIb
ni3rKBbc36wiPPe7URQU+EHWSr3hSJ07O8e8GVX+DJve/0SLC2lBBWvxwGkUeRSpLk9LZbAu1i6c
ox8xbpDD9RyWVM2fbSYM9rV9kUcR+dJt7lb+bVaI9zm52Sy9qq/0fKY2yJK4jhKeO+cA7IywN0x0
qPjTbizrPyf8ZLmjVVc8Gwg2C7/f5QxBngpTx6FFt0olkRZCwConYC5n5GugNNDoPZtNn2Nc6kWF
QnG4OlKLNQeAJvrC1VqNXDK8K3WJlOJ2r/rgCe2eZiFUpea1edcPbPpQdTdQc53ko7wkQa9qpDY+
1L2HZkQRfhQzPmbxbW4AI/iUyl7GxgHiATy2ut+tnRvV+tZTQg80c5e0sPy7nEaNdUzQvlx8QOuO
AnGdYCDoQgwpvi3DGiRmmakD3LdVh9F+GpUpEEoAsshBzaMcHbv0BdutElz017Uh2eIue7PpKMCU
SfS69CFKBp/e/0FHCpWCGfu7ULP6wR08HcEcfiIBu3Su3sJpP2SKsvuh5wzsM9WDWCF5xiUO5bXh
hMIzveOcxVC2Zz/Spr8FOkNU3cWL3Cyg+oTK3Ez90A8hx8FZyeqHtPPniVp1VLiiSxuz5xkEcjHi
eAAyNv4zTsaI+e3x9/IxX2RLAVt8Y6j2T3ffy/hFnRSvoeQRRD4/CETDZKBgDYlQBX1myMs/+nAw
N3Kovn8sV5DOViUYOhkqgIPQ2mv+g1e4fRj5uTFzIXE+yUQ66ifgWgh/++MefJw8TCS6LpE/pWCZ
29wcEaangvIxqaLED72jPWq0094t+cX15doGISu2YhZPyGibS3EBldPS6rxJpbv72hZJZ6I5WTr0
2dmnd8PvlndPVJw3+bMS7eiekQIaAvTYHyF3nWdTVQcSrx0OSjb7dqIHcN5ukC5TxlykBiHLYu0A
M2HjeZQqb592T5xIdpe9rlaGW255xm5FrFs7lZNW1VeO4su+AsK7+sBow+Db3HVv67e3lL3+ozbS
z28x6gwESX0hMqDZe0Qa4NJkf8IJ5TzqPuvGtTPM4IFwKUmxgVWsBh3ah4/BflbpksoT9LhRLKJI
/fwjie4lRhJCX6a9vwPe9vlyKIDMi2VmphtC4sK77HMvqnRU1UVvlbLx467FaaVoEDh2J2lAFi80
9L7RZ6nV+4tyNtK8srp7NHB9UPpBVj0Q4zsk681Dxxa/gLmBV38bALbSzRcTHkPwjYebN4wr4dqk
D5T2rTAV47Dh09oIgYEXugKOXoalBPKKa2WeOXmvX7890LtL973JXMr/7i7J6aEhVnV1DsqsB0tv
LV1B+r2I2ABkhPjOXPwhnozkqgK5+rLsbZEErMAZEfoI2GFjFyCFDOwqcoklxdpp/Rg26H3nmF6c
SXuaPogu7ufludTdhi3Nrigb6BFbx3N8F3WGVhHQxbwfwRab9H/eNqcOX+UdFiDs65wpTWROwGGW
T5QwHaDFSW7gdZWuMHCYuwvNVWuIGrJxM0QEOBcIVnww1zWmwjchL+3hRsm+OZK4x0Ky33IHzgSF
9mNdxjKF6m0Bnl3KzC1cpJmdV1dXwYgSjJeBgDYSeU1KUffi0exlrWrBZBRC3VYbaLhob8GPmYto
xS/WUtzyh06PBBWmILqUOMBFA9xBGd3pYgM48GHh9dbFZIjyDWXXrrYTdfcMDxnPPVOI+QuziTH6
TfzbXJLsqEd7WQcl+fI7+j72XxcdgtvGkckAq7hkLd4To9H+x2dbLkCC3SmPvI/zyUPf2xsq2juZ
Ifidi8t0+U60zpHEvx4nvYYU9bkOm/msSS8BU9L5qaTtbEG//Up/0zl38/n6Bz/Uj5AGUN7nu77n
8qUI1xYhlh3D+UuFrkXdjO08nGMvHU4fH274Mrw2vlvgOA3awmvlSJmIqlVyUdVQMFV/99ZapNPF
3EvO0zd7tBhEM+UIOdIk0oRIr8TDqop3/ybwxxCLm2UCIY3FaBv3z3ZICtBAXt37lzwYNhjODpBQ
Y98QJ3u536EjHnIsfUiJvWqWXXL0bp6CIBIipcGWcnSJ58owxj0pNeyEwepQZpSOHnP0RNcrsuIe
DgxAgrYbjuaFTMxsFX/7/q6DbZ2I1AqZNrXnXq8bNO/5I2YhQeNk+oEl58VMM4waXnumJrAdp0fy
Jn8yp1Xx+GbaBTl6K12JZ+Uaw17pgAumu8i0qX9vgrKqzWXhO7YmXPFq4hKBtr4zQlQTeOqYqoGZ
NrlrHE1FsxsSvjit4g/kj4gWNKkDtg/t3KHJTAl+mBL+l8ECS/rYvdbQTzPW4VhxdN6e8vJ2m6P2
6N9mtL2Cp+eaZEFzS1mY3SMR6i3RSLIz7wF5Y3NTb1WNRx0zr6lI3FBWx46ci0zxbkpHExBapCwa
+6w22yk3Pbn+0ssyj0gNUZTofAHJjn7ARIr0PzrHJqRL+ZqXd54tmggMGvSIQD9eZ4TcwCBMNo07
S+lg75sFq40xAKXf/rVaRdFL/GqhN6PejdV6cGrV2rxKsFDWasyUqwCnj4hWFpOud2Bb7P06Gc45
sENcAqd758V2ke1UM6R2Wqh/bP5npm3JbnRGFdSdJcAkTwLbR7OhOgblsDSfJ59O4hXM8DAzBiRN
99nFkVNi1Ajn1Fth6h0WJA7UivgHw13cVlWgXekfXZQg9J/rDzVrurABLxRoRxyCmbAHOv4kbIFb
YTQ4b4Xs9x17RW7llX9sHVqHyuhclc/RTNTBHqvLkJ6D7MFF5T6zShzret0vC+3gucy01jtoTFy7
aGzZnjAerTi3D559ss0GI1TvEzCS9zZ8DSgmayRcQObm4fdfRtLRJQTvAvYx1Bi7lnDTxLhM8+Kb
bZ6+MeWCOXfb9BPfvFaX2ccHrC1O9TeGrYZqBO0BPNkpQbsLfVwH5HhSKPxMsDXLsIY38S0t059y
v95C/BL4BoivGEB6a00uVZKS964uJUvydDv4NgP4r6EHDeVdEGSu9eElq3vWn01b9ygWBTSWmB7U
OjVeKkMa7jRGeD92lb9sXt1xvFkJQadziiKpC7a4ZDSh3uiyWBpAjRv8KO+0xPhp1tOg3lEOaQMG
+J3OTBI4H92YFqatUUpsKpAq26XQZdyHq4/tBT3DC/UMogi8CMK6t2QmEMQk7JI1tyScy76/mV14
PHCDamLe8BM0ivQTSsFP+KNlGIy9sruKAJqlIaKYU7KLmZ1dVuf03wOfn+hBaHVNXJ2C6YlT8OGD
qWCHFZnXSADwjpd+drgi4/dTmbGQfAcRIqRM4ePoYgKIMP11jFH2qv4RuO2WMys7OEelVz6/GxX3
cRyouqow9cMmeCjm4IvaNcAFwoI11T5MAuTyFZvStQXnvbKXYPtXGKJ7g32xk8lKKDGsWbSV91Ay
Zh52d8NBTPEZW4DJ74vyWesPg18QMKyzerpzLdbG/KrSf0Oqfw8z7bb5hDgMxwSBzLQ27dtJd0UM
qp4OSm2VnTnPXvguLmO8ElS1bIOLtFhfbz8FM7TDLq1K/+COkfRwvUCc4nMS5MX0wp2L5ZxpwXOJ
BwXm413Ri6MzRs+xaCUC+aHVS7q0qG++SD5KTCnKvSKsxv5rRsmPDAL7TKQRWVBJ8ypu55qiwmk/
rjq13Pqo9RskMmdgPOiSZY+5VZoU+vtp7LOHlGTNnYhm12dD3d7I8oONtl4CH9vWRNf/tOLFP7oj
wZXNnjI52vUQqOAFDvu76qk0aky0T5LhJczexSQIVw8ULx7HFbyBVYpMzUR2lgcAB9P5kPb139NM
531a+/llkzPP59k2GN5CcZUAgEOFwxbJc58/kRGyWgzMWHEDiy/hVnc7xLUAr8xzFek8fal4Mger
FwvCdWiWvzuzL8KfLTTXGdXRS0wDaEWshSNoc5THTBdnJnyiFDrPxc1BSSesaU5jIszu3mqe2dnP
UHDVCtuiTfyQHskttFKP/4URObmCCU3qzE57e0J74MNPo8PCHlgX66MOU9FyjdN5pkExhy1yI5aD
i+C/CPN7O5tOPKcQPqsvP5WcgEvXW+GD3eJTLx5haUeohYwVOGCWD2gwmXfgz33SvNN6F1uS9hxe
tmlmmDvTNOuGiEypkKHzoDVGnjWPRjs4iyv3OKdU/twqZSuVbVwPh0v1dOaCQXlWtW4WnOBuKcaH
8uEoZyOL2f5DpmeBiHgQ9OrFznZ30+w14iaAvJeub3TyPO4sL3ueskYlFu0ka+pkQcs0yQP5Zowj
m+rjGh9YCCZLswBEWHvNmGYAJZNYLXjS1vAXII2W7HJSgA/3ipNpKDsD7SUUvN0VPSAcoqnjAIHe
lAhiirp5aNP73+iMZbp241wYTa2SgJyT7tofmPLo/995+CJ64IZ5hFAhjkR1F8jhH4R1eBNFWPox
+z047I8tjupxG8hiriqNfgKMBftzLhVvnlX7A3n/6s/S8Co5MsMrgoETBRhE2Doo+Uarb4+1zl7v
Xq1cJiYr/c3LcZCfME2WZQAfBoHnK6c6gBDl3cblLBgu976iUv/koIOZ84Gqd2zm2w00IYpKkyLB
TAdBFfqhMZjEngxPo/Ewda/cpoMCnF8ZLDNQk5mHKCrKcLVu5riBmpWkbxJEIwGs7EbinUvDFul6
gUcyshNJkfZMqx9B/pQBhOH1jUtTC3EwGXGFvVMQoDmtxv1XLpSzLAVnAZb4GjZlGXf/X7Wzl7QH
nfLxS4t6Cbr/kZw6gDloqxF43sN3X8WqniDX5qj744Jsvm8pxCYN+HqmfZapHFmo9KqdT6ihGFCL
6sgBf/MszGKBdYpBz0G9+VyLC9BUe12ftksW/ntXWE5Qt2b1KPG81X9fiyxfa7sLzn38QVV9jahZ
EY2fmFBEGUfYVSFYD9NF9Txf1PG3qj9D+LP4OoLlhHWHhADlp1AsBUB2jxRwVxRvWX4uD24YdRpm
3+KVBp0/uLpiuv7/xM6MnMrqdfloBCQ/baG51vTsbYOfxoHi2cdKUFa69V97F4AWYeDGgg00d7QH
RkfHaxuM2mZz7J+kSCCjXkKB0Q7z5xNobHFMLLPlZ2n4RauLvChFjhYFJZ6CkDj5D6/85RAoPASk
DbedkwvYHo/mnKwMBsSiPV4D+PqGLEZC53DzzVadboIUOTOXP1Kk/Rk9/812oTBn2AUjUh2ZppBH
mU+Qrd3wdRVZYKcdZw46JPxyIcpc5VuRea3gAyfoDgdQRizt1HiJ1gLsc++wuXxgGoW26M5LMxnT
GdsQ9QgdalQI9QxGR5ZgtYWRpWlFhbEWRhExkjR1Mb29ZRtea6tnZFaO6p2wSQMQK2fsP+eKskGM
36ZwdTJA64VQaOK4yB5ISFjk53oFyaP3TkQMAeHwLCZR3UfNLeinZDTNhmDS+1e4DfClnAOYft/U
0GwHT5TC17tA6bXKPOsKcJ5cwQijh5Hk4Ar7jD81BEak4BRrh22NnXTyLho/x/3NDf4PCsmzLUmo
SuKOlYLknpjfweUaD1jDmvf179feIubRO3ti5T8En3iFZqQJKf2GEEEMI44QLsz3X5NZHSTd4gQk
qnoLgwwyD4VKYv0lOx8G/SAu/zW7Y6oXOOGlqBxIpbV9DhGcNqNAozt0hyehLZcx9T4bnJLgjubY
z+HRhE3GX3OQW/HGAFgxIY0fvrXHpB/xhSx3zcoi2wvmWnx0Kq9rLIMBpviOq9irNSfyrU9H+kt2
Ns1Pznu7ckQeMy/7kemrRzYQfOYhRIoK20dKme+IkUUTUxwYaAowTu8CgbMVzDLh7Ra/uVpZKaBK
1jPzunDuDRb0H0see74mKBUsEtpzXpmKmjp8Jfnr8s7olcjSUZ1TiN+6jwov/qaBrrvQ9z0igjpe
3x8LTp3GwFX0szwKaTz7/4pOM78O6kCVPdaz6dDJinEmDmEogVOKOhe/gci6I5blm/+t4U3s1IQI
zgXhuK7uUWT4dgQWjqG1E3YGjU3vCfUUq28ggRkOtAwy7LuJ6dUiyHpd+ZPHsz6xM4YGrkpQh5GS
N8f3Lptr114uhGrQO0y8AY3eGl/PntnOpB2DdU3zhqWTOq/gvoAcMnEau34Kx2b31MnPEVNNeyrB
K2BfqxUf8Q+uwDiLISUY3gvyUVgOk2ybqf4WLhI0q6s9zT9BvTa3CGozhyHdFoot+olUa3cN26ZB
yzUfoV2VORWWO7c9C+mIFaumRWgJakAeo1rFFK85rvZUpnMuuEA9KiNQNnKVHHMhXpNT6rbX0N9D
msckrvx1Jy0Ut+lWaJjueSAV0XiM5BhOFRCj/WQoAkTqWUUHpoEAxgGd0Jy1bT2gHsFYxwpIOlQP
MizYOmzRlTl+HRDDNL9BQLQL8gbT+bdUFQWjsJyYA4nSCl9Uqu+67s7Xywg35iVVrG0UnHHfz4pA
5tz+IUYVJIHraPi1plfj0yeWQOoxH4Vrl+EYJUDHEFVUEQu6wKx+LCKYEmxaN3W1PwppWle7l+2c
tE6nor+XN8GvD5SYPmTTW03a4xkPY6ypuBW+ZgBX6HPe6otbY/ZmrsEevo4vs4QQ1eG+5vNOOfCL
SPDMkaIfJaUPuRh9uG2NSxyi/OtF2P4KUbGTi/SSGzkfqGQ5acuL02GJoEDRBGELcFi1F4JATju/
ekBub9VHVTCgExuggZa2QaHWxZsfXmdt4ZTra/AOYxouv3vQDvGtTB1oDfhZlVNuvzvbx3bwD2w1
Hi/xW5zikh+PIfuSPNVaLjPAgUQZGsvWZXfgteHWoUY/n3gOXRdXDgTPJ47BhspcyNLpsAXh79r4
8lP3D79bRdQWxs9FQmLKlYL1gi5COkncgLm328g8FSZ7+0cdDg1++vpaK/DI0R90wxwHT+90YPrE
GhcgxLB+P2T2YR72Q8E/MvPynT+MTkbNY1Ep7SMT+yZTdwaYCqa1hRjZm94S5W0UVNvnG3yr11cv
MUMrBySJLS9jQHacRHpQUJrZ9PSZyvKc8z03TsgY+ZXsadT13rQZGMylAxvBBg78b6i0uZxv6L3V
225Bx2r3D2lsCMv4k2emYsmXsFrNmeUHXGHpbGoMkw10LtL11S3dhHmcK6mdBP2zaVVwpIWCR7M2
RVErt0PjlRNzImh0T8MUe6W+mL2UaEq746LyRKcOQEqo8+vMyvl83jBvfaHNOFS6RIltArclZhI0
u50fO0wg+ij53oCANlXxub7mUuNQdHKz5H0p0l7qu6FQPONs770je/jTC4H9F+UqoJtiSL9LSzVB
ALG8jxPCYKj5t9wn6ad9XaJmGCca8XzmUl+EDkU8XuX9yzvPc3gl83eeQC+qS7TL8bH70hWu85aI
mlovAY8toSA98Tpa090yyfPcxbJUBF+v7nz7vYws9bPbdTMAiqoq1YudK/iGzYvkfEx5gPHDAj0D
DydmT8FAM+lIBeWQPDKQB012jRR7LqbaeNYq9vtXUXl0prSC12j4DaEVYMQLdEPxFrnZlUah0oRm
tfwiIl4GWpT7l9LZKADWUwWVcRW2etBBlEBjOfKB1rw+Va2y5dgrqeqsBlQZb5fOMszEKq3zmpxI
JpaUCN0dZVha32mbkPTPCAByozjifvp27wFs/UEXZM/eQJwTkbWVs7gmSwUMQ69FFKV5isBmMi67
TmnyKkw4bznQC7A7hiVgst0J2xIO8A+kwWk1ECjfgZew0t6vluL5axbqngQONABYCNz0238YbBhq
TSFQFhQ3ZCrrk3mnyhit9NN2Gkb+xzNLGV5J2PJFaRTSy//9VYONoDybuvSYV8ikh3bish8iVFeU
2OKnvPIjBmnrJBEAgWjoPup/SbPK44HOVVeysemyuoZrHhjgbgYe42nHA3Ofu0vQNFWpirLMOmUc
115pWF3SZnjeGCve8Rm3LTCdGtY0yZLTstonEx4ivZV9JLMkKkYmCJI/rLYb46YbgtD7UVw/e49B
WtHedavoTCdhLdkdvUoKXzTZEl0iRRxpp3pzw8LnuaW4l9eQaiQMn2M9u/3dvY5tHHsiZhA7h32N
EW6ocPXAaabTmJJ+S54UW183Mt2Ywfa39ihl+5mtaoOnrDoOZM4K/YpizBOsWNKrq3K49wWVRxzX
XdXbrE14QcxGQ+c7JkPLC7VHhIjw+uOevIubTch68uzdfus8b0S5YUVI8HOhI+bFNxN7bhmBPioy
oylZ5/EdQB2bFw1jJo/AKHkIZnZW6wO1aX1tjDvnkU/oZkhDcmEXQsoDRKXVEXsZT/hVZ7b82pTk
eeEw3iUUtKPpSo7vcC4R3Dksva6bAXaC4RkB6nFc0pf4mKImn1wgACUBemTGxsadnRTHpnGCWZkc
QrPf+snVkBE+17N8BNLS14RSM2YPFDZvHkZrb9/z01C292rAxJFg2iuqVLm/88MXEMrGDsO/VM4d
TBjmiX6srOsm3XrJAStvgTU63byf+6v0MFtnvtKuArfmNhtgdgfUo+RNeRWOIEK+ftKFCMW22Czt
sOBLOmmCzePkFaoYOeviWFSz3QMMnDZq9Dj3Ldx9w2TRZzAnGWt1wGVWf4kFmy7l28FEr7OkBiOb
0WFjYJB7SQUTzszzPcXhV8/HWmmPfyvMFInxcBPROQY0b74LmDoYK1P8lFpc08cLXE+sXmyZKMHL
SYm/nBGlT4omosWldN9w+dVQFJQIkz4wtBdvLcob70/352H8XHK87bt+Hg0QmZT2kTqWRnMuW2cb
WG++/36TOCBIq1d2/5eTAsDmRusZu7cKBYPDxTMMfEY1M4Q6zbGKpHIJKdaiRpeFzEo2VgAiXwBc
Z9sixjCgYZttWa17yncmMjPDor3Aiz1a1fBVNHA3rpVei+UqhXUC/4RJ77gjMDfckccFvoskvcQQ
8/34429r+KjckUq6c/y3tKWvkmmg9GoT/9rMFxZBLHElwy0DzH4wRZxVvZ59qeZvHthH7us4XEXe
Urj4NzNsxA5DNeCOceFtA/sUpBgLTAuSKqk1CC88wGhaxIsdecyYgLvpT8pNlQD12Q7e/FgyyqzK
q5rmesAKLF6a/arl3bfDzTSJhoWy7Bu2KttJWWZxSgnSfuALD4dAAifAZUzsmCGBJQGl8QaZ4mLl
3Z3pyijsEW5eTK4XZzVAikCJtWQhjl8P2TBsSK3dm1IiOHKfc1QlKQlrsyHLOc1GxXZ2C5vzXlMr
GTj0bG3aPXbBsqG9FjQN1011iJxHWIrgLbGs72CE0hXLGqRZu1Q4KDuVzUGWmJsYqFfdq3y2FfXg
dWeDK/20ehmZrOdo5foxKNekptx+ELO9WR2r25iDnj1BQFrqv2YV1KTJHp+dcNeDoYNY8ERQs2SD
CFVs9LFpLb+YZcKDvno0jtVreMKHoOjupbAI9BelwEeiYec/4Jq8vC3wKKNiapxbeVp5iwutdQPu
72dZwlGx1rzbrm34M9duH6RexPcd4H5Sl8ovylML7xfe3yIzuTCEdj0e3Bik5iHyZamH9KzngXz8
1XZd95nLjpR8+/r8f+ILgb4gnA13eM3J3W5oVmyST9zFS570aRgS7ZsFAQDqiI9ITSylChJ7iVIW
8V3G7Xa+uhVfgucshJ3nic8I8RRzDeqwJtS8FXvbP9eTJZ+B9vm9Q8xWkcxhB7qbDmDkFXPTzJJ9
wR/dXvm+A5AK/Kyfvkq9z2poiu2q/HhoMWw3sqMoAzXQHOGyCUdboYteOK+BD2SEN8os1jcaN8Da
DMi3lBi9LRqKzWdDJcDmdhfp5XNWGf3o8hb1OsQwoALcGU+BSNik1h/adJeRl5BvAwr27UYiFxVZ
BZXrWYISb6W/+7VWcSVaC49GtMY4Ayoq/+Ee00GLWHh+IPCI8cFdKk3fcxocuqcRcV26mhJIamuw
7P2/DaxerY8J+Xm9HCqrOvuiMVGmvGZu1IsC+7pqybLnWW+WMGlKYUoz6qtJuZ6fCCW2E/xphM2R
dT1Y87Ge5L9EMmNLk/Z5+fcv2x+XTaCATJoCQAOyEbf4qZG687YtJpgwAIQHBWoK8fbOX6wiTmpQ
1rGQXU30Z7w+ZstELbLCyWjI+Oxb4J0emOWLojkXcdIv/ZQQ8deHpB3ry0cdOSUlMA/lnHqcPaTq
YbxVbIB/dz72SUwUqdp7CgLial374RgOUCAtPm+b8VjghbJ1wwEdUVZKugOEA0Ahmb9zddLYrni1
HnKSeloVt6w7fQtRp3YMs6LHLMZejCV2+CH3rDVaa60tgwZ1HjeXsZrbifjfgcbikOjbkdNiUsnN
E3/lAlXlhL2glsjC6Y0Lcr/dVHo52wZPFpSjHCrwxUQjqrp/TCYnIO+tKjfKiefX/ExNSRzS6bnP
NPp7EbsUJUIs3wUTVIiqwbmRn8T8ACuq+bOfylJQV+FeZxppmDLdVSwQRUFtPsEyvjyHyZZ0krDK
+tssinYbZs8NOYbGkbhR57a6UbbCsfTS/xJaF+nnEkFboxhE1NtMHGWD8lzF2r0YVNRagkHLVe+Z
f+r1JlA2D2r4WIIZ78aMWiqOjrn01c8cb7tVWw1OFgq12wf6H32aGcLuA9K35Th9OF6R4/e+DMRV
6pSebvLdwh5NlPH8WAhbBFu3StI8fZLvtyldGoqWO+LYxNle3vIaiKNj0W6INAn/ADSdX/05crmW
dgRL9xf01c6Y3S1qAtmc+xugRhspzeDLczu78krLgH1Hw3fwyJfprdBgwPCg3wUQqlXQRHBsatRX
rkpCo3jXuXH6iHt2ZZvM8T/pfCrX5JFczgbe5RadvTTb0v4rmZSK6aWeNjhHq1863bPZ89yesMq5
xL42h424WOOfpkYo3tOsZB9/Pb7dqFAHaAi2DIcGRtnyONkjsZl6ZLiOXI4C6hoPDZHcz80YbfKH
OxcH/a4AgREkaggr4EtHdzHHkm+kwXip/PidDm4trqruZFpuPzu2KkHVFiwL4vgKpIEPSu+zFGIj
1rst+6TdpmQC6N8Mn9r7PDUZtegL2i1Gzn61/6Bo2+lXVAubiQoYyvOiSMZxE3AbxJsp2xaMBZK/
iGlPIg9iT0TaiPBf1mA8VRKm4ZlvbpGkpSArQNjZjLzetOP7f32ymksHrlHCKCR2WlNFiMZKIcMO
WhXmqQ+F4zPdO8erMJ2NE1b4XteNIQC+5OX9NcEq4cEUnZ+IFAZszUZUrdqZT9M1kqxG9HcaQHcU
57FxRxCDeGpwCwTfaXeSCsbgMZGPkvNcj4r8ZABLZ9V4n/fWNYhk4X3DU49yTWrYL80WtC1I4YxC
c6EP7Yqtz/4M1hN7pAGozBdQG8EDI2QzfzMy7T9aq6bu4bxdICbN9puRPjbOhLEU4lPZSFVk4yiN
L362QAkmNrnJE7EkxSuYpjn0BSF47ml9r2dqb3QaPDt66n+Ruz3JPKCYRL/UFvgbowNrqjI//VaP
uDXHK3sxnrzlo/t5UHDMS77FqP2D8u+JVkCCcXXVpGG0ts5SOVy1SRAFKKAXaYvVr+im1RgL+8Zx
1KxYlxW7zwPb49aZVNh77iE0aj3DOgcLG+e0g6mTAvRuEtt5cNKG2a8ULQJgRF//kOgbL4PjcaO1
D2NoTgV91qQ+qc07cMJQwVPLF9C/jM7Ovmo0I7/HWXe6cxVmLKR6uZAH+fPvvRDvkGbkJ2vi2Ez0
XunSfkcznS0W5CYRR4qsAxx/stW9F6n25I8k3KEWUdh+Tx/XZnQoJ2s2nNz8fp4UWYO9lkd+8ueF
KyMlVjYoG6mj9qcRNtGnRyfQWAs4+NSxEcMBsNAp2sSUp8gS6RSK8mC6LaR6FCmUdX6EIScWQ0RB
CNJFtc9Y0L8+J23Ltd3wgvKMKI2lV93nwn0Hfed8mOtqDeqvUXKEkaVsL+l16zPOS7MakVVFX0sD
s6ewKv2iHcGSRDwxRb3+BT3QMlhvQr1LL98v+VG4QJjvV71PRhvjFPamaptWOkRSXQaystDaZkQE
RSCLNBFp6wVEBB2aByohs+7Ejl6VBUGRqPXp6zu/12rYnEFWFwx5jezorYfXdutBhD6JVivZTLrA
I6wca7lTUJdJjXe1eYpDC0mo1dPyq7CIpHKeYqaeFNoViOv2xw+O7hOzsidiFdKW4BJ8u6HzNKtZ
T/mFG7GKO5NETyUrteIByz/fEElZfsxg2SKRk0LZWDtCm6e1a7aXGsDmYAfLq4/Gg3bCq2OMDgrY
u2mxY6am9J1VSVh+aRwjgXluVk9GEknXetJAWyHnIJeY1OJoodJwhBAYy9KZgYxuFxsoE8NHdHDE
+kaCopUmRARQ7i2q4D0NnnLKoxeYfVLfO5AG92sV0sZ/CjmYfsTVqJ+CCofygXFwbyZQ5MDnLu2M
egeMAG7e1pvdkeB19nEcckXvmtPcagQAADd9bzbrIrAXF2qbEnUT+4jBfP2AYO+WZtwZ8r6b1yWC
PvwLm1DJryIpTYilBIZzwB6wdZXmVRlaeSdFQsFrJ5YS2qbi3byx+tmwjcRI8KqBMwyHR6iSWK1e
sLH0FiqjJqOrnvAobw9H25n1EyJ8uRgq+/7fkD/+t7gAuTniy8qzenQuw1yzJZ89aHMRzUaR3kds
YMQF4Jkh1U0X3cUQjAdW1pEGgqqcKmbdgYeyjTBdVjN/zLoC5rjH5vYmN1Ei0UMygvJ2yzWYbjc0
vOpEuMDylx7XMOHS59r58mahpHcrJThXqjPUBjWcjCOY6rI//SSMQpqDcZaWsv+c2xzg4UgUR/Z4
FgBoPJpYkxVejaBAqmWt0pgouZ1Kz2x6W54NxQt7ZpkEqjwi5gpoPFzu+ONjFHX8Zw8kEohlm0Au
aYUJVSZXPzk9Voyd5C5lHaeF/WJOf4FpjqM6SAe03D3gUplmwtFncTzKLcC+0rTJoXzo8VhtlD79
6Zes5XSjuTNNmfhVvu5XvbWsNv+C/vCUbFjK3RUZL7nOMqkxt62uSv7sFJaIE+Oumwa9YYNDnVal
TuZiSwb5ahsXs3jWrTS0g/Fpeg3PE8su1ryNFZ5MBqWzQP65aoGHtiKb+nzW1d8SI2RrDyTQRlJY
thj4JI4j8zLfZdXVEgqqnGHttRgUCBY1SO4YDXsxBuaM7qfy2cqhZ4wSWdh3BeAdth52gh3JaMvR
qEwMxeXam9m6Cd+t64jd5S3xea+CICspVu5ZWc1St59cO+zr0zc1gL0yBsgdLSzC64KqTKfd0ZMo
S9GJ17grHOCs6xz35a4uGXq2dqfncoeCgbkSUhX6q/AsPcnJRuehnsmbS9xfl9hYbk6ktLa8S1tB
WY0JBLLpFPGvKmxWe9jE89tGbn9hJOqh0uIMFA/37THOF3/GCCyhuNFbMoXhObbnxAcw1r/CLwY2
oKfMN02Xs8tkl9JxHoYStSyA09fDGpi6/ClmD5NOGhonp5idT9sCeqqGDynA5Vn2IIczBXnB7cGi
RcxP5NOP/ks0/fhlkbSeIAt7/Y+AVUZs6EpZZx7rRxCE2ETu++Mc4DIZqOai9DrT57S6DnmBaK1X
mNMB1oVK4lwDy3m0jZOPQK8xGjLNow4mVnzPMnX3YGPF2dH2xyKq4AlARv/9tGhF86LriHZizPct
+yG/6lr54A0XqmgOIdVsptBai2ti29OpBvp8MrT3T/VDJyMdlTZH6gTI/bncdxYuzX1dV45cLvAK
roQnMlgDqUD3re7RXllagX9Gqgstf7PmVFMIBqTXsA81AXwqkWc0Y/Ol2M7y1mXu5dWUL0I7lU/7
veMSo4L1Z/a6EYsZY0imf330gzHE6e3V4eMOXSM7QCOUKQ5vSu2/xmKtO/mVV9iZhhHZ6hVVeTfT
xTTW9UMDEiHcXldQtNR/hzFJFtSlBtiqi1JOXEDBvzKcNq03j6R3lcL1eejYfaFEGMbHXQdMR2SF
rMSEjt7yRwfVoMhVJRlkD74aqkUJTTXtk9DODXAnaJEus+dYc/aEysIt1Vjbzxfn0YDedLhQi9xe
WBpiCvprfFIrh4QI//GqpwNn3TzOh30RThgv9LcXoXx4M9eYqUEo7kmEDuLyu28t//xvcLtRWzfU
PasQnL5Cqe8pSfZG/fudXP9FQUKDTqhaIrqPVcj63Q9JmjgLRZkNyTgfNbCxIBQjL4IqYbKy8Rop
MXo+gahcyMDZAN0AUFr49p/PCXo8PvlIwZMdOj+70w4RENHllzruNrtTnsCpjImf0rNz/jNFjRMX
D7UuNH/yPqyF3PrFUXWQLUnJ0ddMfesVb2FThhfa0Tc7PaRLD3VAWNWBbA39N7gBDlk7Lg7/IrL6
Hdn6LW5F0buNNR8GoQHDw2K5VN9f9cTbKJbYjZAOWCvPLCRvZUHl0tAzPg5YaxSqh/6yaMtsBfPx
ouBvNDd9uocMPf7dEAmoeUnUaz5rHQR39L9e/+0//5dyaU5fyyxR0EmfpEvGABlVrPfIpmivLcGR
xDPkj4fHBxg7ol2G2kK9uybo60Ayn8pFA4AddBjwWoL2HYo93OmN9QGxe5cNPoO8FmsQdvjCWdKj
DjTcTILD7ohvRBBp6Efnv72Ie2L/gwnyk/Cllq+IzmWGmJcbGu8ZFOhKAi6CDJh7x+EhVlZwmWR4
ltTBlW0Y4XXxnbiHGARqMQxW1tdR22N/LWKgSC2nhtWWPQI8eOaneQ9Tq7VKKH5lkI+c0kN/xqG4
PXspjVDhDA8qomg1O4EEFUEB4mhCDtK5qjrsBSOL1XXNUj/FyRMGmU9KkalzYFctdVH60iralle/
1lZt4ThmW2UhWhuwEnA5TakyP+qHz1qKWCjncNAjjt5gOgJjbywEuEIQ+5hXFhWS8vrxhQ5WAAms
/ag4hq62KGx9l3WxYh6QbLZi+ey4JOcjAjKoBWw5kOoBEXpU5R7XAX5TYYRRxq1rnFo45ll2KlZ4
XG4XfWiePzFvtt5BoAkW828aGXM8R4N0SkJ3Xu3JyJ8oEFiNSbJ/oWPeu1io8ZlRgdd1xWqmVGW2
x92QBMwTzrwRokF2T8Q5SLTk6fDYigh0lF626cIDf9RuP9/J+tlqGn+PK8gYaQ74S02jYw7wOw8L
flRsAWAM3lkNHo5ZzhRB8w+pGw8jMx8Q8xKlOpz8iDMgHEHlit/Lu7NXIeSudyl810gA/Dzz+GKL
95Twte3ndZ1N3rnzXcE7f92hYbxSpB9sFSqcYQbvZLONhPKYHE4I6obxjxjHsENWJFd8c3tLyd+U
vX5yp0c6TPnDSOLfU+mVMhOvUevKjtyYuKHZYspDQeYJVgTsfjpD3bFUWvjAZ5lGfwZ2J6b/qDjm
WT4ZpAFmKNCfP4M2mXJ5H8mbGAmSHBuKyHyqbWDfGJh7WI/jGoJfzC2RThZXaTEnRRokKdX7s2TX
0LuZoWJSMNpdKUYe0HSThPKbYKJ/dNUWVancQREdxP2mcCYDPhFaT9P2X9l+CzHa9fpDZjBeK6Bp
Imvt+5ZZC3p/aW3W/6DUOSTnMiEYVKC+3rVBkamDjDgUsjGEUKyBr7vAWfLRQRWJxkMhUhu/6vC5
5coaVDAPMq+jK0RHI1X/8yLhmmRg28goGRX43LLr7Vrh9cuEpKyQ2koNFzDKsiAGke7fqGnfbAGC
f2JYGDIgutql5M7ZNqhs00QTzKAhnNlFdWHWouMfpWvPLeHTAkvM0KHKmmhUUUqCJpS8Yk9MHx7G
B/UMyH+nHa11r5zKvY1qbegveg+5LWGtj88FcitU6ZbUfAzOmjrv3rOfkXQYQiE5sjoRvl+iW9bj
IaSnqhqnlYKJOmXZd2Vxdkz+Ht5eg8cCtcfsoYCDRoqopv+rdCr3t8l4y/k7AdBP3ho0wLCh6WIt
y8w3Lm9zzVCybQToctxA99KWg6d73r9ypDxGjoqCYumUP+t1yYSrRquxWvP6MF+Ksr7UUL4BpBAQ
2hZalIOFYLWjaogpbxo1qz3CmXJUWh9jbeeXGCPPi5RMvLvJrS8uZh6k7us9Blfqrbjd8xYcqSqx
0ZlgF3Chs8SXftzitiWSUzJyW9MRsNK8EfA1dwnFL++Ac1oQSkMTJey0dPkFLO6c0VRjCLK08Frb
+xHt5jXdNMK7I1s7BGL64EU3KD3UdIh5TRyXY0n1JE7CkCMgR6r9+ChIFBBaYUWxTI7KhOWu3B6O
vKouUz9WWKS6PwUpG6NC94lwxf+R6h1h0qx1MoJiAPuNJtGZlm2IuwypAXWnsyZOdS2Dsd4mFiHF
wsCIs3N+FnT+P0zPcnvBmJLREGnRPa5jaU9hGYKtw58ZXxQE7yQN8zwE4A2UqxfprZ1Rl9RnPC8D
VfmNVrVNUrqxMSbHJXmgSXodGGR6jYb+ZYB0KT30FTZvgkWDH9PDHPvsAcJQ55BJF2i5MzJ1XHp8
ZWph9eQwupRyCPDJ897o61RQhGF7s6n/4E3qr/VTuIPbYb6+N4ursR+1SaHwxOeWOvlVMHJ8372l
XwSYry3OP6I6ut8vbCrgmf/xrBm1oLj4vRkvh6/1uP67GQ2b8g6pkNQsA0F1pi02PcSMVIjoIeoX
oOHVhBKFCoWwFEe6O5rO4QZS53rTkak2zOndbFN5bUUrPMnoLdh0A0jVLDBbeDyzfT2EuG6LFSOw
lr1Zt/1SRy8jkG0JCnSt7pVv1uhWgPsxLmEnBf1XHBcU+thf0JBKeiA+780rp7mBYOQOf1PKAuj0
Ep1sZg+STZIun6ZhVeQ9wx0NGy20GxrkZRgDRy3671i3n7CyziWM4ShFtN1eUn0PT0B+oW6cPMZ0
IaJ54epJPFpgICo5XbWVIzRiA8FdI2LyKCOqYzCsOKhgLemVc8w50yljYhV2FWS31YPVN90zOoR4
MFMkdSe3yYy7CDcqM5lQjhyneI/K18Ye4S+6YEGZAFNXiLJbaGVy05zek9ptErhoLAtFJ4fPxUIO
eUj3ZjgQSItFWwTMoPByzNve2dWvbAVZlb5LUsiWFaR9hYChEf3FtOHnlVHkz11+J1sbbfPNMLSH
3hrJHxgyBK1KGfdZhFWlB19UlxyvTu0eEEGfuBTza6LSAy5tWe5BrzLl0QmASPFfmSAf0BbeBJFM
CwgvoMtz51gxbThfo1NcOiGi9Vn3LwJtuuDnQZ4/2Own0GDRW+uYzFU9XoPa9gL/tQtdiq7TM7RR
OgN8IIVo2jiGplnVnnrPg7BnCwjXGYMnH1SxTyUFOsTA2GjnsVjyQbs8Wjos/q1N57NCMZtJuST0
qh99EhIztG0W91DgjzfBV6aU1a/CThOiXckEXXZHkATrqrkENQZsAY/JmSZG1bXv2Wm2ju3o1rvG
MYn/znVir0skYZOlokeeislsr5WDccUUeHX7WjIN6tJO8gQeD0UnucFPWxfssLC5n51OUk+5okmF
tAVEpexGGwXaU+n3idcenJrERjIoFPtT3GoZ5/bmEY9rWZXVNQdhfrwSPmDZZX6VnidulGuDVrcO
R+B1S/r2Rb38/VBZpEL0Nl3qrff/jRlBreKM5ZNPf8Blngn2U+7BVs7DvlIxA8I06Zg0nfgMIeZS
b/aeUktCkvt+fQaWvK3CRw69hJF+PWUkVBt01NkPv3rSRBTaFPyPictPnoEcczWwj4yUjm5pZJgT
oEWGAcmrTlmjUfpYEsoVVmvf4rVX17hHQ9ySMx2DoB3o68MRECHsB+27Hj3ZGiUCbeTihgJdJz5u
nM6j2FIKaiIqQ+WNt825gztaC5MosHyO0M/HSen/LJuIAGDxdTJ4d2cXqdDoQsYRR5eIiyj+Bkp8
lj+qsPTYQwXiuo/q5gLeAk79Vqjnkz4jU0eVjXfIDn9Oh7xzjZhUKo6YU3GEzRLjgtlGFodjnlJb
FPMnnOnOGCZfvICIeWK9/JZbQGTXGdN/x0Kbh8TDYjB2EwqXrYhGj8Wao5sb75qNbOOILihtqp6L
j3ZZjDo70nHHW0hXZWmVu7gDwTxxuDyog9e56L33pk3XBCmxwlKfYUjPPLVzDLZol92zjk4JIrbo
8HcO6WTl6K4VPSN/ieNfoXZDssiFm8wZEPMv7yz9pPGDUYMedmaPUrsTpM/T120h2OzqlCBOSNP8
x/uLFMeO+eok4s2fC4bzIGFH5W+VmkwbdzfUWlPgO9iJF0cZ04hNg0CQZg4J/no91Vro3RQyFI4v
RVKYxMUNW7yDBhTJgAuOpeZW6XEEZHxnsOL+kPxyr6cZie1VXwhFD4Y4UcdVlrjS4131QtZxSLm0
ravZsA9x5lE5zFcmjvCDhThUk3qHLExi3H8ZrUVnXDwYIRCgnvAxnXy22oYpIiKs4LmB9iZSOsRt
XKnmy7PWXbz2wwstqaAmoBPHUpPrBj7UOImGdTuTl6NPyGYMKewukPD1Ekv+3xCszLA9fOL+EVWZ
3ULK19fGTWu35JMqRkxh79qkgcNOfTNS+oG8eixfQ1RstZm0rRv4FD7RbF5WnzOBYII75qzASyKg
AaQ5W8U3AKDKP7Ha/wSHNif0Bx1iwxxbKCWhlJxP+T1PEsY7apvyjiFijAi1wC09h2vIYFMGoASK
iuRyfno2FHtZE2oOPA57pmnTTqfEghhxpEajuLblORbXMttsZDEmSBWFt/wC9DyubAyrjbNFergi
TZMpc9NKZrhZtNTUHdH1wI8LEaJOY6OfJEOVWasd4PloIwX3B8uzlInxxwrse8Ws+4P6L2XlH515
t6seutv5JayVJoE3/MB5F87Uzw8z7fgp7hxQ6VWg5CaFc2Law2S758HswhGNWKh+vUwAWemWJ3la
nYesFfZ2wFaRYhkt58AVbKNYo63FhDR7fTRbsA7u+FHF5hjnLAZWY3JwAzKdp5ui8LDUxns8mAcL
8ATi8hwU8kyJG3VE/tO6zvsoXm4YWLaGdBazVEchlwrNlAdHd0ULuLvrH0Oqsma73i0iSHeJgauD
xTJA0H6nBwD0Ejc3FHkBTXZO/LnvE0Nv67DNQIulsR4bpkgfn5tnwoAtEdPykDFIsgOWCFz247/e
PjzOpbuCrLmSMEzSjiOprjQgStnFszQj3iMyzwE017bAxET3yaP/aWP9Ulfxl89LAb76o3QNh9Hi
Ts4LzqnPzhKjaCRbE8gAXGwOSZ5CivYJ9iGr8JjUZLlZBVYF2/pXfJKPqQ22RcvsM2CKdxBcwTn1
UM9P98le6QHW88sQpCMV44o8A12n3a9mhUa1sWFsMIQGB4cozfkr4JUdxpEc6uFiKjCDjsoAReEF
BepgBYc404NRomf09LqkOjPJT6TDvKu+eLAN53Z8F1y0oZNTH0pnGPSqh8/xSsqJTCM39v+U4eO9
ssO9qpGW+aK79sFNGGOFMcOmLuRPOt8lG5rKYL7KqNt+7ONMjBDhE93E84quFnNb7zdFSgE/0R8V
/1G+pPXS63qUfw7DRYztaB1ji8PooPYw9Ms416TkzOMO9ftfN1/7oPn28pKxUyPs1BFv3re0KBzP
LY77uF8H+uQaeRZvQEjUJdZ7bkeMGMWqQa+FDVlcLQ0aTeixadBdOJlm4iqjrB2aDiHpQOriF6UR
5XhXaA2Rrp0sG6+c7tAHbIVWt8Y9poBrtbCZGPky9qX9mPclzCx85yc/UDPxYfk9ta2CzRk1feDn
giKjfDcevQfVuVgKZeXoWoAHAYAURdo/nXuXR5rqPFlqOH3n6Nv2lRO9OnlMoLZjYm3KEc0zGsbQ
9fRYgF7aenE2upelPqT/CJPWXfatMWNLL+YfBKFg9hx6Gmk+Wtugx2Ke8ozcigs1ooc8s/YJkj8B
zbaB54zJXmn6Upo+XKtncEdcJBmPeCPeCYvJeub6amuPgI9WiZMp6dYeqvFohjoeBltR9WOZsPpm
Uu1ai+8Qg0iv0nxI3SFWuOcjoX9dyG3IbuMFmPKWCMinvQy4msg1AeM7ClDKp+FvhtwyMHvLVRlK
XRUIODjyud+DjHybNvBZt4pm9pfedUOyueh7nZucWOupW3ao7EZ57CXFSoCk2kx5EBlqEWdlZ5YP
EvS5m+vW2AZ9zeKW9rVdBYt/A+9o54g1l+zNDmjAg17s1OVQqkKLj+3WUqPJPKKpZaPBb/5HLE2s
xx5i7v91M9cTTINAtRJLadMzn6JFX7qQ8zTL+S8NY9U6nBchIHnZL1gKcYmHBsRYL2Oio/v+vaur
JCDiiYGoj+vYkblMN+StyGJkMIsIf8L0HYpeetuinbV2stUElmaHz21P/NLt5bXh3LG2n9S0b7Qw
rh0f6f8xeZqOZ3f3rV5yDyjH90v5/wGXQv07UEyaAtTMD1NK6/bBgVR3AdXSh0xkZDA/ZJzf9zLw
kX7DDDy0vQJgrjqqA83RvhxsExDMIoknhNrxWpxHUktFk95yMmjWDUxoLwC2AyYg4lb87440Fdvx
LbtOiMpkkaT4jGuExOqFEP9oQlqzUGY70II9gpYym5SMRDk0AYGYipTa/tYnQYoATh3a7ac/ipi3
6YlbIcZ1iKsmpDoDqeYzMBiSJ/dZ/0o/izo+JxSznWCcvPD2t0jTsn14uNlj20dWuuUSCoiqh/CV
t6aq+L5DI8MBf68O97f2Z2mikCM8mBIPFZ2HsZcYH0d0CqIqG0o4YnPVnBVr8HV/DP62FWv8Ac4G
c4YLBg95jSdXgOaQyhgQUc86miWH5bHVt0NZ/u3/N6WIBcs3L7BhQQ+cw2IvcbNhMG5N837NT+k7
TSnq8BdPidre6gMRYrON45n18Wr+LNbW6mxLA1/J7JcxNt5PV1PQEzI/edv/5elmf2ArtX3l70uq
6RATTBNft3sCanZTGsDPZt+2q4dhBQ3EHoikz5rerj+g3PBgC80AsRdIu3Q5HJd9fEPMLC1IP4LX
Ayee4OndIcWyiPKowv/laLMGnfNv+TqakuGb2Zk5PJfKXDUMjDqFXp/OCUTsDCa7dl9OY44zGPdr
ZOAjSbtHlIWERnK0Aob2TPLl6CJsmOHBHKK8JPAjaU0zwVjawh40y7wph0pcQyv4Bh+jP/e5AHZw
ySOcakduw/j5xZhO59flv8Xxjt5Uy/pwUy5K0ORyV7hkOwASl3AiGRDZ85F95BtRQmARSjMDAlYI
5DqjBWohJVcLTu7sremQGsQacV9+ouPDOLF3NR3uip2xA7lCRTS8+ukW6Fje/eDwflOAmG9axfAw
+pLbrl34IJYqjIjR9e0sL4aqMsoZcaKoqCqb9JSJhEke7e++YybNBwq2YZJvSDqCcsm9+neZHIfo
gqjJV3fEfGhZlfQLMsx2blVAA/nrmxAsMia7NlsU9K1xhGjOf9B153rXb9PQD+e50RrIPESksK+H
XfIE1azpkqj54lRUvhZamTbJj4B4mlmMbvytLMhT5DdvJqLhZJn0tGpftqM8scCmmAoj4Ir19z8B
THeisMw2L6O5+bV5l1LiAUYkIZaIBDpvQ8kIB1eH3t0lDOGHlF+gsyb0W/ZWkn3QS+0vjQC2HRIp
fu7ULIeWkzNYQPGD5ZaFdKZTFwDkGBMF6xv7FY+6O2D7jEdH8bpoSH1SUnUOV3QwKSkBGPsHF1vn
wzp+Y4SqFP7DVEVo0FiG6MwXYp/nAOilXsVtOWvALHSbUq/Eq/T93qYd9eRBdfDiK7soUMTScAqy
YishbeN4eDixlGUC5qrbEYYUejYwD40CQH5lHRjF4tUWalDRdujHkZy7nLYkd//r9Amunp8FerAj
4E3KCMdQNMZzDRjyNMPk/zRaxOS6C21BmsWmH6JjIDUE7OKGjaoR7qTgqtugnCJeHU1mxjrEaQxV
658a+q1fmoye6ozrreHrgB8yhrLyTDzs6LCaG+PlXjIwphAhv2POjESIXRMq+diFK+I3gKKeKQM2
GRsDZu8SP1+16foJmURlxhHArPDa/KAPCYvqNB2SI8Lkhpr19I68SvnA584UcPWg7H1rnDWBcHIC
wHWYL/wf7FmJ34wxU6jpNFFs4Lx/1XDfgK3zD5x77vjUzQcl4BN5zhOBeVF2xiS3gn33wMnryUa1
JrFruXMeZtniBk2UlEtEb+20wjv/91IcgE8Na+u9U9GVfSItkxtPG1BpvPA8QFPgxdvMikjIv9kC
0LZ/wWhMJ180R50q+QJ4JMss2rNqvy1ps7VSg0QPaX35yKTws5rnJCHY1LZV8EETz8IXsiI9tDA2
n9TxEGFYK8vYp5kqmgNDKrM8h6dtMex8wauM7s6cyMWfjduEGQnAPraupztnTqHXHRAgsDGC9/Wu
eMsXpBfV2VgVfN+lsoGpoMtuJbkWO5YNQhMU78XfQo8yCm+gRiN4zVkMtQC9h5XmsA/GzsoA8r8M
BuCRddatceWspTUTElYWZqCjip4ArX7gTgj2Lfdra8DTsiBxuH65McqOjdnxbibMVLjTY874wBdo
vuIazXNy7b2ScGN382PIMUrvhd6ty96kjIEEe5pnWTeamA3sN8t4sgnHDbrXBAfcaXpxqx7teUb+
LoM3pDmVNN43jBkLBMe3oSoCG2v3aqy9YLSVhsPH8lTI0DfQ6WGc5ebAndDxm+2xrORDKJE/4anQ
OTdcsGPq+7iEbaM3nF5g8O+SzgmzX/pa1bDIWX8S3ZHKN7mhqZCyJH9AjrpDMpbhDyCxBQqZUGf3
5YkdUgaI8FcM4gxh+Eg/60PT6wO9MwsoAPQaRWIMcuwIL0IZPcRM+yk570Qsy8E+pGSSXstpBFKT
Ya/k8HG46id7CgOpIeiFSQteZpGlDgAi0EWVhuIGqPDwXYoMT+ga1E/ixUu6eqHJAXBvgY1/gqUl
5Bls46Ee9bH/pKGadpLutM0IRohvDCgRtyCla/hKj0jCdp2YPl7KI+KVtMQAoiyWw2dCKuNBTQHp
BGTV5LcczHkLcBd/2I83cQdZnEUp6ny24ihRNep7U20nI0HrDrTduo5hMQpXaW3r3S/t55fZcVxS
XulmWld7P2NuYWjkxwDjhRZVjy8KAQFLhjrU0ltjKOV5ubbQCCoY+zBTb2iLD7RvkODtfN/yrtdv
aso47+l45TxjPIVvJZ8VSAjz1DTH5BR35NWUDMCvleaPDJM/FlyL/ZmYKmnIRDv07d0o6TKVOwyG
57YHUHng6yiyO7gs+tGU9I7DdAFDzYMLsgQhuuk/MELjUGRiBMhZ1FBz5MnCQeoAtL700Quj5tyJ
9MR78oLQewv16TEOx7Guofr9BiXTTCZCH4e2EJQcA2U+N+Tu9IN1a6OxONtPxYweBxsrLebw1Z4g
Y57PptXwaCHg323xc+miSQzk2a9hDoKis1qA/JXhjTtEhLhrWS45j8k0nkLsPzzcim1csshjOWJC
12HMo0UjQY4FKokcTGbZPOwpfDKcOBToSdUhyFivXnttE86/C6T+lidMkTXh6CL+ZvmE4zQOYKHo
hIbgo+vOuOjxOUY7tOc3JrbCylaWsHDoUQg7TfF/F9W7KeIHfXsGRXY+4IUj76umygKMF+K5FJ1n
YoRNBXWn8QVCNvyoLnDSs+RftsSVg7VSzrKVDHtOK8XLVVWmyn1X3rDQS/f43kMBNRuO1osRU33k
8WU7YQ72Ld2RCo4OarLyHAPEXi7SPuiTVYGFnBy0MSgX+zZto1iVEjE7Us80vMwKLYVPghg6Dd16
kwb184c4HWXwXc9fqjj0tjg5MWRc7G3tnnDSAa8puQMIG6bFlAdYkj0l2b/DOF2qPPQiz1EAz70J
5xQ05fNNnrVvp7LD50RyUqD+9ZncWiI8blE/OEkkvcBLcgA0VHP6Pl5PAQiVGFkBPxNyODTZ16W1
s2bDduYTFrEClhNjFGTtrMmGSqJqVp+5MB0TMIaPo8Q8CcmINVyuc8zlc1cnTL7rf9BiFwaBLLS0
QXUbuj/ejCg8m3GGCSOMNK8O8cT5Q0hSC72JsJQYL8IZ7NfswBxoAlpGc1Je0UcLAKmeNTg9/uKR
uOAxMmkR1J6gnFkbGNq+GC+nUJIGoD4dRR0FWAHBHMjhRpvsO3vJBmBVaqPr0PTj6/vQj75xHYJa
g9vugfwWOKl0iwFnnRgomhtyAtS3nEOVDqpnT7pndtGhNRr75cEX/73TYjbehiixlLVWDvtwUihs
+o/n2gDfFoXvkeLnrnNG1fKzJSkyIZrjpUgvQyJ+r13pe4L5cSFdnJoPqTIuf2Pluk1wVYgTV0wC
xp9YirVr1lmhRhZiICdX1VCjzrQHaFu3HLT1x9hvVSXA+CElCKC0qbgLhz2KjHomstvVOYFsr35e
XavcVwgdcfEkUQWqHTYyvqSIjI+bIEF5ZaWH/KHT+58Va1zMtmvncha19CQ3hPVlXoNlKSxCsVSb
dfm8qDRnrZh6WFts1rCu4G5PcOi6tQEzOLkOdk6x2xCKndQnctfwucub0i9ctRlPckcwjgSk660Q
uDnfWMwTRomft3GQzZK6LGe23KhMuX7G3VZz9YrLT635qgOiApaSIcnLRBDxesm7AGUKuj8va3Pv
Nk6EU1B8ODXec2O+Hi0mf7A0GFdyBYjsitfQ+DltXykBFu4p/8XXKIDAeLqhZTiMv1tybl5cUQ2E
Fx2kDmZOrQQz9GM/QqWyaG5TAMSwOXXrD49wjkhEp5uHOZOZMhfn/GYpcgfBJJo9aioqZRVj0Wtl
SPwL7J16Eq5qsK64tRcxFQ6ormZyjlrVU8O5AsHrSN+BFtcbp7BL5IH1XJmd+rQGJHWMgycYZLfu
5PzjIzlRzRzFEWuMEyqkmr42jkrddADFpsOdzziXQuSwE2RnD7wfj9CfbTamuYP1XkmO16jekc6k
0QPiNzWO7VEGGt0NwNfN2GrPf0yaE27we8aitutNCHUwu0AQ8dyRoHlNCV5aBR6o8ntXtuh2Wmkj
dkSvc9pxbz8WMUHABKrtNssoTHJ8Dg6422jcI6OjWQF2VPZ4HQ01iFaz5nfX+vXTz1js5mgLOzGE
Kdq3EL7vuHm9oDmN592DV+ZE1Tf7t2WxLcsGz6bxoVj2JaAE4adKFSVBJiVrCbz9jesbhkDri2rf
RxhuOhUWtVih7l3VNDTIUrjdzujXHF+mSj8akCH+oSWkc82gnhy9u9tGuz0efAoVfe7gAVkhxF5Z
7ea96WbpEWN1wZznuaLhTWPuQeL1HpEIcAtXsMkoeiMmQP0N37WHX0F7H3h9VAlVBX76yFto98xo
6QO46pf5WD3YcQv9ACr/iH5p8brZU8adJT6l4TjCiGGY8CaOnbZjft2Dl6D7W/rlhg5gDovryi4J
rQUZ90ZiLXGykeI8lUgh3uk0YoiQTWefpI4N9y1DBWgjDmvrRzIdlZIDhNSfgOTQRqFeBiEF3fiy
Ni0iLvT1OKUwbLe6EqqZEJvQOhZiFC3EZ3mv02UnPZf4DaSaynSBydikPsJ7I0E0JXf9jf59N+W3
Rv8+1hgiB1LAV2u2cv1ge7IIeCN4Y1ZhA5hMXprGIeaRHlLgYe6+o0u1dDgGXdEYNF9YtzyUpv35
kBiI19yFZ1JsdYVe2tWHgnqm2fid5dp6hy8NFM+0eL1/bGbyjg1sokk8OkZ8zzPypkk6AWf7Fo76
AQEoiui4tOY+C/XRUhr7ToyVjRZGJs+GHdxl6Q7kcfyy0PjxCk9AmtBF+GRCqyeNLqCnxW5rqQfF
3VTVYST7kSvp7GYwAC/nv8UKaL0A79VHU8+iYI9tGyk/5WHbc6H6lX+F+xDDN3yMTpVjWAnYOR1D
z+Iy10OQtB7H7nSKeN6E4Rd4BLYA/0AVXQ0qgYnw/vvRwTLZ+mh8QmZ301UDOQ3+VvOzSfFGh9k4
9M5mAaFQQB2sokz9z65rtnZDDZ4dVAOmh+JOgZH5TBfvmXbvmGvzeMi8+ev0vxP491LOJ4CopzYM
KxVL3yQiwROtQ79PovXBL3DsdK2XJUvJN9WPf9Jj7+UyJtf+d7IoWciTQzJjiipRtxBWsB+NfwnI
pLIgc2bvEGrGBkj2VaETg7He9K4PRogbBNcf6WIYLhmapx+1q22uZMIQPw4qn9svzAtgyLbFIy/w
WXj2wElyN4UyZEGgHp+K6WscXsdJjuhhh+B0Kn+AEfDfbK1NXRi6t/kr/POxZVcP1QDdAy3wvTJz
IKCkVBPg82+XBg/Y8B5DgLhx+iSLllWHtDrlaCEcr4E6G9Q9GqAcztUYJEaRvt4Cc7nH9TMErcbn
gMQlpUCLdDy39ckT0jEGiAsn68uRDNu+7W3udIGkIC3YN6aGgU1lUNt9lpXvrpXUKONkHizjxxIH
vQmrK2ZN/OmtQAd93kzbwt8liPMmoS8cdMErz7xz50L981xQXonhwLlj2/L+5f6oWN9ml2irIFaZ
wtyG7qm74qNbBQjiQgFDgTj3nDdUmhp2vXfFejj8BBITyAi3wTHcCiGJgnUSdY+1RqRhdT8NRcW5
7GeSGOqg17V0fdnO+j2mcMD0vK27ryjXEscVopMisCvOR8MtSNvkEGOzMwspqqmcEt2Wi+KlrvIh
gh+TohwgHynxNENBvBDkEzYSKx/D1OFnMiSdSLmtFvASe54Na6KrrSoA82QD/0HS9R5UawEEiWZ1
1xQLJt8PYQJuO34SgF85DjSQM8+59ub+1Wt8LNaCMnoYTM3uDRj7JhovZ5SI+p39MuiBJWOF86pW
PRShjfJZvGQO1TQOe6tEyX+/34XCqtvS2OTXVm/N3mSulxTLL9LNVpLN+HM+iCJW/ob9UJ2RcITV
lnk/twMgbf5DTZUCbBEciRiSI3FUOLSraIeLb7YyF1nAA1hcU0kBGCQv0FMleU9Igo75OI53xQRO
bcp7m3jG97h52qBGMurcRdFXEHBZInt0RS1fIbOur1Qjnlg45UdKPiTSBc3/V0GmF/3HF2QcD/gv
sfPD45IdEsWKSNj+YA8/ACwnodAKM01ooAcedcdQWfl/UGx5bB7p7HDRHxI1vO6YKbMRgNAtWz0m
FTazG3DsMsVZT0xnMYSSwYLofSDnZR1lnWQ5uv5oJxyPUKKSlHW3kQTBvNRh6WYC8yxHE6IbVOA9
fqVkEVRjxA0hwc5jPOr6m/T76rT3vHyYt2JvlYQ9DvAh7D4xNSyXa8aKfWiF8DF6w61U+q4yLy1A
v60WdWOwq/9UsuIVaosqUls77Lc0vZtG/ImJu+ARowIpG2aUPcXGQltis90z1Iww9Bcgb15OVwkf
4RrH313VjlAZ/O2k30zjeiEVMKHFydH87GEMLyXs8YFrpGlgqzasL4NhH+U5E+A01Apm3Ch3Kzu6
Ix3JvkPyJ8GvCZH3XCjOY8W5zG8/LFZQOUPOba/y2/ZR2lpdA9NwUL7Y2k6PzezhQef1mMJnXtxX
S6Ym7dCLACfnGGmf/hpZkDfCUkyZBYA62FWIxDe9/k54VRO+BJJP+tObQrQlrOl01qO0VxKUJTJA
QZRKMw01YOJjJnB1pMMl9YYcsbbMt8ZkyknPwIBlKqCgSiqVJTO+lpXQwiQBEcy/p5gLHk2rKRmA
gImos3CkBtviIDFOStyeHVei69Bb8bsN7OnA3jE8rbQdXcX/E4MEcQLzVwPDGYEb2zQIPG0cqhEE
23KXvcY2WlrQl2/PstdrlxHVWSTWtebxj08UhaqaW3B10m43qWrLNesUUtZSDWd82LrgHIJDMJQh
eKuNo9XVDjOL4gIJopzIENcugLJhzLeIrCdTV29146VNVM4g7ZQhNAgz1Pz+/R8kqla0MpRiA+h5
4Oxgpqui9Ihdhh+Q99di/g+MTyJ5+yLKBrswfiqabwc8WUfBMYgB1uoRrRQY99yZELf2rFH5ETYg
NZ/HJHt7pfyzLJOwSg3JqP9r0iPpnt2hCtB0h13rN65E/Odwje3JC3fVfrmwsu0INkdA7GbdAK8N
gZrWys8oRb05aKHw1jMJwfDcW1tyjRV0JcVPQ+dAuybdJQQYyNk8AaocUgH9MUFL25zXyn+WX3yW
6iW2HX9mj7PU5a8o7aKOzgjXiaTprkGBgPd2wyffk7LFsSm6w/D4ZT1BFwwENN2LmkAQRRwD8dte
6abK+dG2byqfLjUuWNBcdpYF9Li+unVwfZgYDv7Hia3IOo9rJOayLuMXafWohTSuBAKmC08djdlc
AOYq9lYkwGEa/yP7JxUXek023vZBotkKJoXito0x9BA9At57FKIB7XxXZW39SuZn7YJFRhvBxUot
niVAr3/5GaJpuNvm6glLLl3BeYlr5zIcaB7cGXpF1nT1OiDB3VAoCRiR8KdJf9FS/LRJlTcBylbQ
HyK3UOSaiFuL5n2I0PbmjdoLnpeu/yku2SVgaZTSiddYYW+jHH6ekA9P2MFnY2JHiXBtfkzBOEG1
QmIqJCM5bWYfSP8h4tkYKVou2ooWijBnaEBy2uribCuy9ErMJXmTncgiqN52+GNMZiT+g0XykCrY
OMW8bLXyw7EeHBY2r9plEgRsoCIWmZILxqownA2Io/Vl0gbqIvq2DA5LO7KE0uPFRJ2QN4C/wcCv
Awuh50uIS6gtT6w9T1RF+15Xp1JYE/wXoHxmtL3jUVnkf51PrySE60N3MFRt6B7Zk/SEj4rkLDOV
MdtQnp24agRLkRrHYXiA4Kp5C9jMkJ0lr2SnV7/oVn7WTasbaHj2w321lbaT8dy+lzw3ErSQYacg
gUZGdMkiE1oEdlCIEnbyYMhetk9RhEoixxyfYz6o8+6m+2JVR4UWPE0ni8BsXybYPs6Eu/4xAvDE
ae9/2WAmzkMbIbT9+zECV7S/XIksWAW/7Neyowm7om5Qdx1ifJ7nIEEE0ky9P/fT6S6HvgowM3rB
TUo+18lIJ1BNzu0ftDW8r8VkLopEFVGbHyFX6xBK1LnQllBQq1TUmd/BtB9wWvTQCuINgE4I3yxo
rCkI53VoGPv8mYgZOAlK8YiQpN0stZhs5yMpvW8DMsdyv2cYPfzanja5ZvM3xQJs0hdFaiTRpH++
ezt+9fYx6fUzD41wWQU6UIO3uULm9d0mdt4iIC/tUPs6xulRpHwTOLB5kGC8hXmwg/ENa6r5S/XI
7EUEDBGA0EVZkZvudAg6CP5vuuQuhsXxP0Lp+GZC+XlYTq/a2GYT1idQsTKxqv88aaQZpg9pBsqn
ec4pqdRxtxIJ9jAHqa7WkUqcMq7OGOyt/eLz8GrhlLKK9CqJdvb+nJhSP58x336k/Ke41ZwhA8pE
Awp4OKFfqZXFdexVtR0jbluRm/vSjxmN3sLq1c8aHmdi6lxxwscpE54ywVnz5BcgrxILLWmTMwGL
ibF/wVQ4eORBh9d5Iamw5TJHU/CE80yDebpsdMVhPljc6gJiiaZseVorul5SAWlkZg69ImrKgADG
FXpKJzyCB3XVGYKI4X4CyfUcLF7eFpNPOZ9BYfuIitCioouacI7gpYZ6ZexrR53U7BucCtVOzFHO
Z0sYpO6N388yAkIEbchyn0qtFJQH6Ua9kx4ixJ4UAACgXrGFTEzRpFqBDp33KtYJZbB2NkSH7f9c
W/UiaARfVpDthZVegO2b1NWss3IfGhJzspvV6UO5bKXuKVGNBV9G3i+tvngLejwZ0qMAbT6ahsgF
n3H2EGLOiAiaMlM0YVtVEoOodUoyRv8v6FIA3eq0bZqq7wWmIJJweixip8cR4ajzOGV6YZyP/hHa
jqnthmaTwRUx93w/idvpPqt5uGag1Pdgj03EHj4r6auZhN12xI0kSxfINUGJODOPtCmKipGWcWw6
0U8VvYNlrkI758a+XzygjfFav1klkMKrjPNMnrRWXbcW4Orv6UmNIqlKznk7WxhghB+5M3MRhm5a
Sh/r/I8kRlX9uaw42uKL0jV6BQHMZSw4S7Wfac2rnSPRnBKc0Yegeg6mnxQtK4LkXyoDfnvXwXyB
rb3mkRiFtk7+z2PvJWvOH6ZQ3zezDKygxyGhuW0ZTb+/iqbk2MHr5rMC5dH059iRJ//mle6wcQxw
n5k/+D1kySWKybnKhtllUZyfOnH+TI48eRKqXKEkkKLtN3e+ZfFBMOWWKHYZEXCNUKGaK2AwBZSu
XDZJcGAJxHgXJ7zhG6QU+B4BmobjDnAZRh+5oA6d6Kdp47M9QL+uUw30Fqlle2hvs+V4vnJ/dOeM
rhNn7JR4QUjpnORH7UO7YMQvEt+eoUJG3OqzA1zjGpOE6Lvsb7i8BdewKqYiwJTpcRwmPRukFQ6T
e69ta7aaEJab4BsmxzRe5NgYmhdFrV93fhSshFccmRp0LHXi/NOPeSQth49y9IUAygNrconE/kZd
EGpixXF6MxuRLJ7OBhmw0BBtRVMglFg+Rn1/cG6cZQ9MgdTfxSzl4ZbVZ2sz2hDhuv7EKq1UksNv
q1XdgHb8YIy2ZL85d9QYYVIddK7U9a3HdflArqc4cOQ2re4unSUCAeaNP93oyf8XS6Ufj0FAHcDg
lQlFE2fH7AFSSrch8oV6Ur8xW5cQHF0zWAlo0aWD/NVWU8JsfzDAqVnz2729aGUHKsri11vfm67E
GnF3BR5Er93Fe0pQNgkbXYHGl3iOSV5+jfpXCTkrcrAHYb18A1jHIDaFJW6B2cYjb/JqPvRGFdm/
+/Alq3jih4K5MoQ5RwOQmhSo5ivTZndCs+kmUD15AWdI/SX/ubOCVC1ES03rXGVYGNQ9fIkKwjY9
FBe1VfSlv3MRrw28TedgkexmLf5TW2d6UQz4BNTHttO5UegTafQ9lvxsiuzXhEZ/pw9CbwYNZTgS
RDfqVIGRaDBmveaHO+E/0tcnj7nI1LzQxQzeeNQ8cnv8+pkyPUCK9q0uQQbY1YQLlxaDXRvlXxDc
m+JzHSEtQkrf5OQ29l31Xq/orcxAo8HBsAwoycmy2+R2IwRtfJVCrPhF6O6opib/CrtTU/fN1C1d
GEGlZsU6Fa3al0D8M4kf46zC364izrGm245PzxwKQPyf0z7oLIc6RHYr0qnBjUCfOqJKL3Nqm9q1
kiaCzQ/8kQOQu0rP3apuW8q2DO3C/lvNjXLJBiMYBVACzzHwIbQrzz09BTEh8xXOql6Fh29vgmJz
SwJTK8Nn3YwzZclYTonNBh/c/J+5B0IVQ+2kAGFkKEdYt0coE7jnR3iy/E7XSho+F74C9aSm/Wuk
pcWetts15DTLmI4F3ho6PbZK32TR9HsBiq4RoFu5y7cuffZD45h1kzLa8Gs0yVZdfRFOS/lXgc0V
H71JLIbexVXdTZG/MMLkNMRVBmoX1G0cl8GaJwpTHtgyRU2XGVLOKqe6DoKkwyyWKLvPVOG+azz9
SjDW3qMGT5Zy0vL9HroiTf5w0bD1wPQTChJaCoyNDHY5d9NtQiR/OkZPGh0VAaEPaNobOY8tLeFl
5T4ZPWf4mSb2TmME++nkFKRAZR3MkPAgTpMu1EcTNEQtcdqgmvb/Tg+Ch8UGIqty7YOBhNImJbH+
4+COP1yv9EUvyRzdGyMpka3O4tN+3QL4uFCwEVWY7A07UzwKiOmFjhIKtj9FEVPmSJ2wPVgoJapF
hBPtSPaupH2XljDwtZC+Ovstvk+bCzn9wJv1QexJb25Dhe8p2HpGeSvTxJSMD8a87VXG70PLaUZC
d0ZhDLTVGZcl0o8vO/vY4mkwJAv29MKx3n2InCpDoyws/DwfMCx9eSqY6C3lNhsqWlDozSv+v4pr
FiyInJ21chcW5ZIXmIIpU5M0rcUzChUwYlg+naVsmHHyfQtfSmRruzYQqim9G3MceK2ws+fMU2vm
/qLL5U1a575L5gFWpY0MzwTNS+nSC3s/f/Acu5eWdC0BKA3zl7bU1RUOIwExTHI9BsK7nCEKX/AZ
rjHr9pJhJJIUQbgVigJX3/lF6llAwLnA7z9df8UMMFTbiCzqd/W5RRxJpIKXAvCapCwL/QsUDZow
LaA5JsN/4HcpPsIHMAJeXxIXaCmd2jZI99idIlo0/pe/GmKvrfIjPHT0p+n0kwm2KAcmfdNjozXn
yooemwTqV7PJb4Dq+jicTCedeHyX1YrapOXkQihqkKBfct3mU6O6vrQO0N5YurUrNXxTvl3rOYDD
uU1a7IFF5Yx2nu8uTdtDvKYe+oXmoBcfNNhNWkgqwnNVO+jn8S8DLTC54t+PmKgCKFBUsJK3XBi4
LFD5o8N8YIZY0JUfK1KqECuujePjFe+Loc5rbp8C92/PABVSzSog5WFpE8dzz1JSCDqTLVtFAGDH
9IKvzYXzbuof8Q7JW5BLWcmbvjgohYmnaTEQSCe2iQpu2lsS7sYvs8mvEf3rGy5Aj1qPPTeWao2k
goOexgHf5jAHf3QOs10pVZpKg7nx1Ugj9OYSOYuIBTRaaUtSxqwwpWD37SRd/NHyct+zMdlL/AjS
byW2YdfEZMyjleXW7WXcsBhQEbN5WeHbslrzKfHI0aH+wogw5k74ULr77Ac8UHgi5nWz/jGPvCB5
PNw3ZBvKJhGsFgfddWELo9r1+Jw5/5JR37/37t/DENcCj2rtG9KWtQ5q94YVIZU51k38yuz9P71b
/4TMRAJFdM2eyugj54/eBDVQgeno9jFv1F94rJoDtzUH8Breke6i6dZJUU5FzwA5z7OM+rLx0uFi
hi4bDUIvBfT2OHzfCTe7oZRx9yAildr0I7wZD8Uqf8gymJNidAjmkB37tsjrXISu0fax+gL8y/cl
3uZ12SlPcwkyP3O0efGHYVLrUbDujm59jbT/bOWMqXt0xqAwBjMZ9oheB5kxw84axUVCJIX5+4Uq
FHffJ5G8g2CPWt0MC2eUZOGwaAT5ggeySUp/65fZ62wzV6fU5Rh6NUazPsrPrnhkyQtY2NyyAH9c
INDNQfCWg5DHNsWkVu7aSLIVPuaceNZnVuNz+zw0WKnyxvvfOwCHMIhOd6Zacp22sUFih7ZO4M3B
drCgVnZR0YrA8+Ufrm0NojzWRlSAG/M0gnnO+Q//q2dqFshrVeSgltrjoc1oG+6x4Aoy6qaL8tiT
QfxOKYxwntX8bL4XMc4BjldBoyvnCwhM3lCt3HtcSyR/xHY+xgieK38uATkQ8FfW0Bgd6x0BhgiD
5bAHHvRgV9spKps1cljCeemJSrnfhsdsDrKgOZRosLLTgwZgnqXVaI7NlQL9gcxrshwl1SnzuykD
Jx3no9tCRlQAKovGOIHQjFLRgaEeEE6qddsZc/ELASDIzc/zvJsCO19rXc1BBDK8WQtgxuuk2duj
forhcOyySxkTRGBqdhdrexAbO4umR2XGFNuur3jaPGynBdWRND4n+7ZS/X8+WkwkrZbZ5PUISu1R
Ax7VuSkELDmkrdtSz+sOXZvtLWJnLvy3MQNMxo3xszc91pAK2xOwv2L7tuWynRgEQ1lyJIIpMRkS
TcIxm2RAysK+GnWeYUlrrPGwvM7FAJoUBI2CWxopFiHRy6nu29VEmYChyNFVxh+KJu6xUAr20VwD
XjSI+tDrWcKyiG0GdX+1izixQLbRmMfUdTSlYJc34sFi6qXMZTJgasbcy7otbylg2PIrJmmtKgL0
9KJ9jYXWluQcOGhmM25EYluYb9MEwhJmKMKVgohKSurYUOXqZjiAsSSqgXlsM5s1FGicgZchTdDZ
0JIEOIXUXbFyVLiRLcXlPaxeYBpGPFzTEu6dihoiESS5bt6mEskhSSxOjO6fDxIdv5jRvijV1Xk2
qXnoT/U+z1L5w0lOws09it69j9BJ0rOr/Mnu6Y61bkGnNn2cS2adpuEeGqTQBV0Fm1p8mFws0txu
8GezSivxv7v7HK75Vkfm4PHV/Sjb90I0IUb+yf+IvbDCcMaz1fD9iUZPdJPX1OyqRoXJW4FeeXb9
Sc5lh/NtT57f878UUdfw0EHClubFlSYG3RS9bPfXbblAyqJRxPSXoUYkbkAM0CBz3Xgu3hpSOt5I
yGufMcPUkuYUlsRZAekbDXPAEJ9NP9eVhT1WwhSrdHdtp615S2QR+1aBK2oFKpVbIGld9+pC6HX4
0IXPg6QTaa1CaNhIszkDhJ2XzR9DNHVPM/qhihuBvWIZjz4fxpWOvMHHO+yhdPpTmS4TMcdq/Otl
B591FdaeH8zGpRI4P/xNbiUOGVpUNsN5+xCcBrYRBVrVckcpG488ulP9xbEd9kvc5fqKIvNAGyBk
sLY66J0WHi8xvBbm0CXoMAmRjtmUQAReaWaiyo1PTI27PDhNotJYNnxypBHEhvLmkC9YTG1CgcZu
cA9fuKm0bwczBbdW1ziTh15rJS5bn5YUdegTTqY0yVGN7uPmXE8dYCc2o9uHOakmCdVI4DM5szUZ
7d0q2GmbuhbA8D3DfbkX+70HdqFrkiZAVxtIzjcgo0N1Chch4s7v0wZyxXoswWQRX+GVxQ8OwU+O
+dYWj8dsnhJwhJz6bhXEhch8ABlaqckMRfUKtgWi2Q4Nfu3zJuMA9//mUuo4aPc/kxkZjmxp4SoE
S7yuA0BOerGdjJLakTrOkf1lytTE+q3yl0G23AJiXmFXt3lahen93rD11N5EIau3UlfSiuBJOF1m
n1R7BRMZpaiLOfVP/5aoWh5zvDLkGdpb0lZpKWBHV1OAbzSOFCgRazQ7xSUVIcQPDdBdrYF5GXg5
zk9v+WbPMI/YCxZJpFBR0uP0CjR2A5UaWcQ70xpXfSy9EOH+mks7blo5xi8ZNsWKO9iI7UiFBHCJ
KfH5459K6ROC4R/3AaZ0JRiyJxn49NtoBn1rpbh1Sgx//xPJcTVEUgJE3FPF6Ql0B7BtEXKHEQ2D
0j8XW4fb/G8Z5TcQnXNbmed2QsQFKXB4KOAhNJw2TLkWd7Ii/U1b4o4Zo/8VZ1v5xRTwoY9mDcIa
B2UlpaZR9GbsiLeSc8uZfVJmKlVBwFIUhWLBtUr6rXfPJnViB3euIMaCjNyar9GqjcV2fP8o3whA
UdU8HVDeKazvCyUT4agYQPPQiTglZE9lWMziEYFQoi74D3q5oug0e6m9SJ4kAuUBQ5PPLe/Dwt9r
lc53N4pk00xF9suNk5Evg4Z2FUwvX1cNBm3r+X7KY4ArB1xofsoWXwnKime03rTIkjfR6L2+5ynH
z9GdTs/h/dVNBOQWcFLfhpVwtsRwOcws3hdvKTuob3x9VC1ycxBQ923oWjx3BBRIgZcEpPhSpI78
47G17D+ZbB5+iXlBbR3pCimi0n/dvN9xLUniJVrKuiXwOhCBefKqdL4OKqaQPrDtBnUtfv/x5MqT
GsWh/njmvposUWppJ3UeX2jHLmgdvph6JmGxOp7J93rQyF1sqC1xJ56+sIP1v+hpKoHNIVZMk9tD
3kUDstwhnXyr/i5xMjt8Jm5Sqf9qiy/NNk6800iJBvq8R41KWQqO8MQOZgFgI8ZuNfsHBBsTHu1T
D6umGcnACexJSVITipCQPUoeUzEbeEmK5Be8QIE/Lav23Wot4pnoxT0TYpjSPVVn7Vxzu67Arp/I
OByxPAZaH7h9zomwHktYNv8ZPzkeHenarhabYdx8t/UdGvKhMPn0FinXGo47rJX+BHhwRVakLNcg
8Hxsxp3g0Scq54fBaqGC7H4y5OFbeAeYYeEYa7VvY7mmNwcZwlgfByLUciQ04nacbxTmDveI6F4V
NFrgalY4kijQjGobM7/M/5gJ8kS7er0nl/XAB0778SMjCIMhLj6EJdJzPnueALhzKk7gNq9AnBAi
S1aqN5CGiLBmbkZUlfR3K0e8Uo8foZPtFHGKKoAIKIHz+HyfPBsfrDcL500a0f8W1hnBD5u6w5pB
ButIWRuncUH9bGspmEwbIMLanW+q67SguYMRw2RIJLKwDJgqnq7Ps8UNLDsu/1VWGhXRERuqPEUB
8a45zj4JrKgoHjK86ffB4l4Q7Tg39v0UBCPLdoRpRLDz0bj2zuEcX0xibKDHgUt9lWOL6ND979DM
pHkkDEOJ2gfOeVExTa9gyh/rWmjzC1NyLKBeSDa0NV1Q4SmZWiGOctRASDHIHt485xefyprc/hTv
0QiHaeFs2TyVBblZW4SW8HEjPHc4iVWkQvPHWoaQwq5dJaV69DzdqQZg5WHpH5Pr2tdsVDff44Fp
JvUITgFpxVg0TZCPS/gmt61mW8ngrHdPJnULajOiTrzuB571NyjRXx15qtBDobQGbPMisCWoTXEH
p43+cqx6sccaDayV+v9bXsAYZRHBTHVra/DkCGQAYeeNqGJzcVfzj9bpRdbIye0sWLjWkna7BOPv
lDk9kqIlJvKL0PNv7qMGhlyrLtFRn4sm/2yowZeUqHQ/su83xLNz3x7VNV5kT9t+5WyB9y4UvqbS
f5F16GoRJ4CmOzhEVn7ZXheiyPH826MxdngkoWRZTnVPIFGsBsdoS9RY1GydC7bXJdVq50W4i+vi
1sVqMotCPPui9GXDiYugDSsd04lqHuaOAY9OuUBxUjaSCknNpBttKhfGCpP/NIVAnE915oE/OjwC
fSd+BRk3NM97MNpaqU4hqJC5+N2T6S5GK8TGLK1S9hXGNPnQVPo+qPRAVnzHTkClb5xMgDr7tTSJ
tCJTQ2Xq9oS0f5yZ6/ky8grH4i5w7eZYGP7goxEnEMiDTX3Prr8qb55i3mLaU8GIrt+s8V3By9LK
qvrQ3L0sJbBAPEjh6LSXvR1Ot58u8jDCDYf9FSzIO/U7ZJotLj/J5xyI1erIgKIJNPSmh2GVmydh
CfN0SSg0mC7x7rY3He4azES2bdHAV3lWqrDVn9RR1jQKzlm3CPC+CtIbsi2itSvDTnTuu2NmDd9g
Sy3sBzdCuRZeoJEaCFB/UdZTM/+owHgxpaJt1JNtgMi0kSAKMlUK3fxAJ4JjreFVs9lyHjrqutu1
UhZDWPb1LgdXSeXFflNxov4l44JFfy1szjoy+XI4zBLT7nspDPozPTpdrU1sXIXXxoRvB3J17EFM
bod7tJJiA36QwSDLfHcj15Cebh+eaMAf9rcZDRPMau+LT4Xw5+n4lZHO5LNLhmlgr+B54+IV3Fmg
DQ30CTMNc8EfxvQr7PTkJ1heaIV3p/PPUInysUpMoZvLGjFg1a1mJbIy5M4l7WeoazEhAPPwI3P1
r1awRJ6ZqoHhZ4dWrTdcChfmZvoqO4kRdS/QO/W7EVfqO5KKn47oU+bMTclwF9Tvknut26PQA4Hz
Mkfc86oAiYz7rnJZopg5zQyBGiOhk63tBpycm4fBdoSllQAPsX8tube2aKkBPLVDeAvUftm5j0zT
oGJT3w2DibS9ci2S5hefGpLq3Dcvf1o14yngslvN78AOJE7bHq6/3eiFbvcfiEAl75PQUs9IGjDJ
ZqlFWLzSaLuxru8AOcFvuNTpQsbUa9sIEN3roBbL9dami+H6AVVRUfpULPV7xOWIsJ2v8Fr9Hldq
z23iAg+p58mSrsdtgfV6CsxskhzfQFuqiOkvO2VRlGa9Pjz5hrRYEfUbn8YWzFvvzi78xKHVTCrd
IrDQaSjtVGZU6tmwZavrCzmm7mFEsM1+FmfgOEVbQGK/nkFZUuCw3rbdTI9vNiuDSQ2/uix4w4jj
ySGXOo6cXQ1gjnIyR+VgNBoLzpTn/2/TZEyMn7Y+FeuBbmmi9w43ezYeQspgiVECzPBjO69sU9H6
jl5VxVPo2rCmak8Y79dJbu9chByhTa4FUCjqLJkirNpKp0zFrpciOYj9r8ZoaXuWuJX8CYYLhyBb
uHVgh1Fwt9KC3JKn94sDZLcNhHoJ7EEcZE17vrSHyQ7Rbteuli4Byk4YFCPEASwZmge6D/V4eB7C
9jB0HAcbIKjpoYnVMQBPDNzm64QcVpKsFeq7KHuzoJxsCkQB+9pgShIOPKnWYllnrcDrNLkoEzLi
7bfNz3WNqcK7EClWnb26afGz3mhCm0xVhAs2IwC2WxBZq6DJ9Ue+FAa2Q0xZgu4YboBlwPNxaBJX
DA1wuMftgGxdWIAOjwNVcdq3kG2VX7BqHwSM1km5CqyrWvepiH6DTqberLowZivmOFUgJJU1rNVa
yaB/p1RGlWczoY0OR1BGKWiKlmeDkPLXMUSdkvZRSFYSkm3O77D419XS63nnJw5mdnQxwG9QxhSN
rEik3SqaO+JafdkAHc5mgZpPGLpE6k2IJp9+JeftgT0RPNPTMfowoEdHAt+17ugTvsAgYAHMJkZX
tLvjo2zoTVI7kMQaIW8qFA02XoBIfam+K5c728pRzN6PKBDwB7keyWMo0lZalWFSaIe31gKvO3ma
ibYTUgAC4xCKH38SM2CImN2v+XX4WFPZZOQKjlDuRW8YBSN+IFleLTJoKfrKNRGRg2MKWnyi/zpl
ySBqxiUaMIahjsfl0V3LAqpJ4X3XTquL8yxxxRo6CBMV2YHvwFXhDRTcqtmdOvYiKQIDs1l48skW
DIVHHuV/iyMMpTHqqnTebIZPQTTg8k8fHmSDvzR7rZR30cN00VsNZPB3MHyKde5PV9Qx2jtVKnnl
o6BgEWf7sSwhgdffHqBKZqE7jlGBs/cnk1/cgm0kliBYq5jVkro3s6fFGmeI/AbH026nMWUpwwCH
eh1/VGPP0SKxlTC/P6oyrLUbCLoZ7Mb2bv7vxaQZlsk4IjUH1qe2IIy2wqcnhTmn+8sEduLR0Ym+
GBX5k6d6rsFWFM5CHpcMiAhOL7E5srtsX4Mb2gHQ8PJra7BTaPrDg6ThLrgEp/QYjwllP7xarUDq
ENakfNUvfFKijZBR6fe96Sjk01AERCBnh7W72aHNXP23dHpV3F393d9pa9Q5xqaxz2Fxum4fmCKw
1XJMkOF5/3IEYwEf5bCHlzr319LAL7cAPxM/QQ4VJqVzASzeeqVfLuo/nX3mhzHnuveFw6QkaYeV
eCRWbEHg08qF/AoeUDt0rqxrfSdkrD6wABczvjCK8R4OK7JFaMTSpNX4wwsfc2JOfa9xGHdy3JiY
PIcaV5fXkGFJPfTHE00sfCHgPkPeas99WQb3YJ/LnpukN8KcU6s6Zxa6IPdsDjeKyxqJTAPq1HyA
rX52ePXqoZ8J51D7n4kXH+rPPBfX+9TuY14OQuz60jZm36eRW4QP+tQxLnU51/VtIK4VmlRpsqaL
YLZmna2TGLUrY6colFPx/VCOU0dhxWi4v/xNGIqhfBGt1PwJhQBVb1CQ7ehDzvd2fZcnz8+OfvLk
J5nQ2dyONuPKus6umvL2VikTAFTInJ5Y3gptAPQV5C9tjVb+x3oNF+HiV7rwJAE0aajW1DGglQHB
DKHphglLSRe0VSqTVkEMbnNknY5kdrimlBxDzeAprUEPsF1W5BMEgSNT6QseSuGOoaArnJ3v35QM
hAqOkOXvR4ISdEmBw/BVRvlwPBTulbbS9OCjhj/jdiEtZBlw+aDq6edIbTe5pQm58KIshzFr1Fy9
oqt258jy9HTb946QF0mSRlGe1Zb4g+zD+6Lx1DB4n8CrMN/AWLqIw/GNGxq86NRGxIUm4CgMIzxj
PAUKyFJ1ZaDrHBg5CFBWzr8YvBtN4tyIEntXz/tt9C/333cJ2F4eNbCE3gaZEyhcjnVz685sBYhj
nxir6u5yicTyx3S4ljmzQDxd7+6CWW/W5Oex7yjSseG61ZZmqVa2e+cBS6PshJvbaAJpJpWrlByg
MV9THQACiun9cbKD1tzyu6zTuAzDd7fTpVqD/sqfA0NADnweRH8gfmmtNfVN83hQmkkiTm9v5fKw
W4Ruom2ZK26bdd4ALhCgYz+KVuY7Ibnqu6QqWsa0ITF2sYyKtgHnFyU0t/fqJ+ICHs2C/bIkq2aD
pw7h3hUFDJkQi/WchkBM4j8Li6xKevnxYlxfysMevAlrnoZz5op+SWN+KZ5jNdO5pR+UbV3Yjuxj
et347Dpgv/BO675ufv00BtspniX85xImSr4rE6kJkQ7H29ZPG7BvY/urGcxfrKDeWmtFtczd/WZj
pGv1ecFTrbHLWF45QTwl/nbG1+7NVr5FpDRn9GspD7h/7D0XnrMPkvJJcmnk2SV7aOiD1ffsQW5O
QaQ/j6Nbz9nP2ww7VIGjk7aeqmmPsFLSPMzo2cSVCbb3YIbpwssIk6E/3a8OfxIfGSYQPC2CuNk+
ZqKdx7olwFMyYsjmr3ji3ITpQLL5MmcAfxwmraXEqrfXGG64felKJbb8j/3LEDuOhf8rR9U5dv8t
DdEyLzoi8CHOKZEVm2WYQRQ2HtSV2jt4cBWuafyWZm6s+QMXzAkV6J9Et83f3s6IJd4BI7CTSg9e
/BWs7BVcnN4p/EVUxkyxm00HhfAtUX97SZ8LLfO848NjssydpKeipCtIifMKo5LMzPcxShgWrcrF
A4EQwrvE9z1dQnoEG//umRBV+Uekrb6g7Crwv7YyjhRFh59JWEpeyJe8jKsEcOg4C4cYqoS+7gNw
lvDUUK/YvqOBmT+Es4ZASCessx05pU1cVAk1H6t2WL9XNT97BSxgj4OxrhwcCzZTkfQ5j3uouCgC
q9MjlB1meFP0PcnLJWf1DcLtOZ8gB4FNXyICwLWcNKuO5NvhWUM1Xyj5ffzwFZoidSYg63QxFYIy
/dHfSJ2UrliMFreu1nb9/W/lWUsSaBAJbHR8i9dpRWa78h2KjviO3KA01YDYuXAAVxXXdsMLLGvJ
xsDwwmOsT4avbSHF9GyS7nptjLwjBnhZBoqr6yDSsEJtqfdLYPkJaKEXCJlkAie5IZeBu5ldzsTQ
0kyBV8cCw7ZBevjCuzM0BAbI69RiP0YrhvcA0LvFSaLNShL7azwMhsot/8OJaDplsulYM5XAIXtX
D8WWc96JZBAnfg5JobJF3FPZK4Z4FxIdnYkjuisoXqM3r8lCtK9tiPfxs01509/rxDLTfna9FBTe
Jv3bTh0ApVeiO/LbHFFGq/GsG5Cten1MsxkT+HtNnDPEf8OSw5ppk071wYKNbmafpE1tUq8t1FzZ
i1xCVs++A7/++jpIDKNGMQqYvul3ue+oozs9s2mqxl9EO/IJg6ll0DdiKuKUJeoLZkevmhzYd26v
ZDPYmdjDbzxY5xnveLFAEHr4lj49GW2Y0Ms6deKHnLTVf4BwY6gCRVwMk7kNQkSZXjmf9dpz2+Ez
47IVlVvOs4/xw40IrH9EtiJNu8K4j7sskrLGpKpLh9u5Cfp7P4Nw4eDBudx+M+6L3qNaXrMjFQhb
ZfthnYdTEYFH4fiYpWpw/LNPpJHFpeM+wSfwEnR/GlOHxRjSwfduL9MeYzKx9cuEsJMzIPRZZi4/
A+yRqRJJl7MVOM1iqGsiuYql0e8RCjTZA8RUkCfQt88Po2mxkRklBNO65sP08s3lyOgNV/OOabYs
3kmgMhlhj0eSkZNktFdC5dqOBa4hfTfKvxKBcVrSegSPXK3fkaE3fLTeVXRTrRnKv13ACBVwyg8/
XT5ncfjJcNzxBhXSFQCBQZGI6QI5hjW2uxbddvNydgfIvB3bKSDZEYJnLSa3/d2EYBD4PyQWuNIt
TswmVDxqUB6JXThdWj3W/XQzq3zSgGGWZxB6ZUsIESyhGDv6kDG8Vu5sMHJl8YEsDjbGgCP/U4Lv
Gj5mxM9u3pOKywrlmbbi610kHixNO6vehNANWBV49ivuVAZ5fidUSC3YYlo1t/KX5KWDFJEVlQus
FufEJumP4ijmziHCWMe3cjZ64v8Rn4IGFZNNstDnLeAdNk75pXhzqy6gI1ylhy80KvXglKHgggV3
EbgavbW3jUrk5qhE7IT5av9oLviaDAjlQV3ctA3Yw6AFIZREik9A2v4/t2WMwJGUiUX6pA3O+UKQ
d2P1qU1na4A8jr6cCKM/T/02OupyOg4JZ+h0Yb3Atb/yIwJ+PjgV2K865hAWN+AWi7tUgwdlBHDH
I4j75zXTvL3YQnPQJNJwIEeIqNhY2d69ZmLC7VooWRZyMXwomGhge6YFR5oT0oet5htxFaBXsE/K
4g6mUm2amJeGHqm7uyVIYjX0b01youRQ8DyUOjp65+dZ2eYfYXq4CsduIRdVnZFYOAiE13JwPgFI
S9nqxLetf/nX7xrW2gkWgj9qfzHzxkrD0ZiiiGYTZ/GdsDubUMJw2WdfPMJ2c4WA4jLEkxHNZQha
ewHFQNrBBukjCQgsOefckVD1PfIcp2K8sUtQooLbLijOmui6/33Jq5bkoSv8n2O7Tp+gtkIZCEr1
5Z414ahZSdoEMVzlhQXpIHW8ceV8PLx1Qs1VaNPm6Sue5+ZpuBn6Km5TSsXbcpvuqTblwy5JNjhC
TqSHLQOOU/T6n/3NlBQk/5+TVyMq3c5FJtAwnptXxKg/JMrnUuuqLQIs80Yl4Gms5u+OHDzEJbG/
/WgO84jr9yHKYAb3pI8u8+vBfSt4SUNnB2C7tq6T6h0wLUGU3weLzdWoDNJP9JStQPggEcb4+EjO
EMZP40APLSRHYS7rWKa4lhrzIk2bvJ3fZ7601jCS5ilJa+ZWcR/51tqoJ+8gerGOE/J/ApaJIbL5
FEijLVo57DBsx/Gozc5+/xW6D3w7tnn+1eoHrrkmJJXFADccBXExp4KS3kDtXeDsbB66/smugIgf
MztbZFfnrPDNwrjZoYjEyJ4lL18Fokz1I3pVPVeq6YKAAciKxdCMPMyrTZLpVV3VZb8BWeS0tBnE
90oeI8ouXRLhfyy480nkFQrLKRkHyPBJm1JdCR/EyEOmeX1S9gH5y/1fpkR16KrLUkwb6aARUsbK
olcBwVf4u7Fjd/c9rCLfA7Ld5QAvNLf+YtYinKD8CJqhreDqYa+RPgTLHlS8PgqPnlZHg/MTpUXA
+kYXevqO3fo8jq5h5gkqb0ungqXZnKuDoYhEziczMWy3vG456pQqYN74OVV3KR3KD5dztgXgzDDH
gTjfV0XCT+hBrjvC6iakygHjs0Hc/7q48CxSAiP8ovf3XSXcRlXcEGqApttlCzcA6kLNIQBSD/Bx
AOVXAIKtDHZvACzySypTYFlAAn5q9oe2GFCmW6dDvQEzfdP5lt7X8LMvrpASTQoTAVpoIDJZRzZA
KdqEplyJoXoG/RnPT/3eI41391OkVcT2BCfkBqBks5+jfQDfjwgrr38m7Ym2kj9xhfR4DrGsqGjw
msuhRn31puaiQKm7FAbgnu77hdNxHsmFp72hZ0VGVer1xmQlpjSlGWexW4+rVgB+WoZ+rIk//CSf
BUMG5xltVnG4PhqHU1F8tZJb2s8gxm/pcyAwZEqJoQJX8OLQNIIh3+pzvaXntdDivD4tMWrIrVIu
GeTwuNvgcM11NgVdubBgnDvxmIe7q1ntkIf96tLIyYRODpqcz5WV03TMp93n2EvhXZn/6MxZ547q
hpqW+wtgFbx3s8aMifccktSkEm2DQ89PHtcfFbkRWRZ0IoYrVobHg/39EnhTdlBjeVOyLF84wgfF
Avt9D+SPC06INapZnMYNzZp1ydk5CgTxVc62qz1D+rktCAxm8/01mD0MjsP6you+uio+H8ci0qre
AeRRA0v9y1w8wcjrf+lwjyWxGGkpwhgiD41OXSstNYqXAyJYZDWVqZdkPzd7O6wkZdLDBupmQfwb
wa4+FkP71YdCKPKS0efUP8Fodo29y9NweLJ17ellqaGJSG0pCKactUnDSWINjWKwc6eeHH5z8Rl7
mZUxtTx8GMK5y9bloJaod+24S6vry3R0gSDc9v3+T1bIu1y5//0rauO44Gih/1y0JVDwD7RPkUq3
/bvP+bNmTif1aHSTu07AZ2XvJaiFnpgTrl2NAwa27B1XXhYj8f0DawaXKnA9jd7uvqnzDi8stsz6
CUw+1WS96SWVJ5OuQ31ttQgjDXNd+X80aHyEHMLzqobbwOv60AMRJkgdyuay7P3aDjnH+uvr6WH3
AUd9YOI2E002XOzTbtbvtPVVHDOOh5rkLnL6UbKePSJSlKnK+JZPGv2z/XtL8cQIy56JH6JjjkzX
SAV01CPzFjiHfW2VpM3eN2NdqmeezDT1wD5/lur6Td0o60tXT5VJnB+El90QSmXmevBgmGXtf8dh
hS5E3PUqawDyex3bUPfaHysMgtJ/4x1qEilKHHl7yp4/ZPXsrLeb7IDuEi3Gi5OQC6A/1JGXlFM/
7I38YHsQcdAaF62rUok9PY+yd/03dxAKCtMq3S7cEiIqmlGzOfNmko9OJ1PJF2bhsxsBeHmf0dhG
P7xZZbWlmiP2TaKJjzbvl+JjCglPTYv7OwoyoBUbwtaw6YPrn6YyxUrv1ckn9J2L1JoPUbgztPJ+
pBaZzJG86xkPrG3uHv1oRv3k44cU0LKLWAgrmzp8vexp2Tb0KbWoeLFaRjgxOK6ym9m1M51cmVwD
rwNBnzsp9ZjltpNwEk3eIitQqRe6IAHE+MdG2v/R1YaiwwbSSntrCuRntDwZnMA2l1TcKPaQpsgK
Chb7fx1W5L8+9eIxIA8/zsE97Q142xzSL39US0awBAFZD25pMnaDDhfEgxB7so0WUtkYJu1/lHsg
vhUBv5HpLFO22T+DIHpbERYndNvJGoO1bWy6KoKvg8F5Do6XlK1Y66CgJOFlrXik+Q0dXGWF1PzI
2lADr1JBSwl/miAltCbVh9vnih4ASjEfB+O8oPGVvjZaNwhdEc4Ey387jCl1h2rtZ6YJ1275Mtmm
lTEz7KpXVabxhkf1gtKXKCqJ4L0xqDi66qswN7s/JGdhsVjo0TnO7hoou2iE2JgNkG6ukywaKLMY
JO5jRE3XScKe/mUardQAWjajUZljimWCiLKfciUPMfuoLCU1FIq2xgXUnRnD1QEJOqxAztw6Zlla
pB6719zk5t/3noLEyV7QccL43mWng2F/EpBooPbNLSPUWX84ELpz8S7LG4mkpexQHkJMaeVcrL8b
Q8+2jpR5pPIKAchZ3DlHcpYTapX9emco13xOEAaSdpx1sORLWBIsl+BJA3oQrqeafYbl5lJvvy9e
xHsSDBJPf9jQ/yAtHemva/g0UtmTovF2w57uRC1fZguwVKZ0sYBFWhh8UHl6BvD1YyKcI9Jx/G/z
qj3x/qfgSm71gEPEH5itpyJF4lxH9yomT/OYHORpIx223cFGW7AUXdKT+wn29U8FaKu4g+qKgwvQ
kpGR7HjPY+fhYQcLHqmSEh3wDRTTQsThNWwTEXrbC8Eaiya8mlnObcaNTRR2lCh1ixgd75qqj4NL
vC66BWcJiOSErKej9ZUcL6G/OsogrVplUGarFfFECOOK3/62RChNOtUCYeB45d7xhnkTa31B5hQu
O8k9qPLZFQ6GHpGzdqidxG/I8njzt+dFqy4g+Tvo/skO7VWdvWPBpY82X5HSlE8xHcqpkqNxZG1R
M7js3hxBwiwzxfUuaHjnzcUf4Cps2GL4NbyM6DWUkvOjFzA6CS+vMnMUWHQvoWBF7VoK55iPdZiZ
xmjF+bzPfQYBIrRD6pzcQ112z95E8a5pLTZyhrSm0JEVJVqfIln+hsQQ76PqfjvoNgJeFQ6odR6g
+kr0h4RsPSwfQ/r/yKglop5uWtSqQvf2BQ76xpaVuRSbQggjhGSr2yFc8gKPhupOEigwD+/0NaML
jITx+0wCCXva39wqb48D+7zMraGn0GAoXjAdKwRnqzn3fpyAKHnaG6gAIOE+4kZK0zE/U4GyhtoN
XY9W283rDW4KQCfqicHcEkM74TOGcHDabkrimXmcKLjklhTVW/D3jkNAErv0P6i/SiQa3Aq8PIwG
SHIYq+O1t0mMz6CKLmzXRgEGHWp0QaKLLPUSiJP/QNeA5zQvDCnhF1Go+urW6XUwf4OEPCY9Ksh3
GkuO0iLhloNNg0F9wFyV3vzlpwBNk6+F4CC5eBqmpkSes3MBacaZCI0cOk74KRxnQk+MDR6HLwW0
z8ibUAJEYnGOikt7uygKr0GxublT54/85TmRp++HRjBDof1c515gim2jDykW9a5lKdTGvCicjlj+
n9PRxMUeSG8GnPDxTG/8EDcafYOAbDPFArsmIIDODT4GqTxdN19TUDBUKjlv4cvYtC7gV8J32ucx
q8AG9S4K4NR7aZlYa/sqIz4zH4xPBWZ1zQ5whhzusulGv3BvkGHCWOVqJ0FVCTzx2yeSsaJCD9Zj
p6oxMEveF30aKFAyKnzugG5Bx3mkjdUQKczp5Cx20PgDCI9Xh914e/SkcOa6e/wcxfzML0EI7dzG
2ctoDcRNypR4jrJkfS+yssg88/N4dO6CJw90OTl88rbGk1JUCSX1/Yzm9oD01VjMOYgrquPGryeC
XDUUdqOz7K+DsYSLRDbRQ9kKCxUOYjZ/e3LNX212nZFuU69ktvMwS6wbrZQcmDnyIeoH8LgkH6dv
CW9LVQs0X0fvlbTv/tNucWz/8GKwKwVY2bqHiLCzoJeIAbUqrLT7PRdSbBTuU2Odi3Mvev1NfxjR
NcDE5J4Ng8DTFw3VNmcBv05EXjrGAoDQ6dO1t9Opo0b6RPHG+dXTqvjBQgkwIEAPybbGm0U0Dm8A
mcs6J24rsaIutBujIRBqv8wv56y09efSMOQmrdNyYXl1wWbhyW+rts7tgYscOvHqSCeYODzZhbMs
GzVGvGfUdQtkbw08lll0I8wGqHSCI6lWlHxA716AxTZA8Aj/6aUpNU4Jp68sRDaYGGcjh4lj8gfz
KG2RKT0z4bVv38B+gnD0wICJgc7fDu7pWlLL9GSJPWmefIKjClTuyltXtaawPZfM9F7GiRNkyVHp
3o92iGdiDW6vCNhWt3BRlZj74IkLtDExXZUOMJ/UfF4gDEUYNknfOUPNSkUXMOKlb1KCFYFTLZqX
fGLp+Z8XDgLX1aZSbMoyuSAUheDO7TnKnUL8uOOjAEoZCvvOMX+P21847kx/1pu6Oo7ZOf1amfwD
7YAmxrpftc5IZLhLPK9a740LeXEakA0e8l+yfb7JuUzz8dni2Tu9tis0uwmdYopaWPP0xtZ1VGxo
SQUH4F1qAnq45Ua91XwHifm86B8cEBqUDtTkasYNpDR2tONXsmO1yMTxHBeS37KTwOYgnS/bZOhD
Mm76QOINnCUSsgOkJ4fKLzfwEX23kr+3mdhcgaRcFDOaOJQYLTfyhrX1VqVQHvEaW9y0XGgGEmya
e+EzyufWwdvizp1L45rx2eUtPto+BP/StCUWkRyDVewshd2m927wOs8xy1tWwLNCUF7OHZ73M70X
ONtDjG74HX8xsQ1aSqFnMZQSrpwKPosDU6Q7gYZ2cyfZ2fXPpYSk10lbgYBK3tmMytvc+7OM87V7
fZceexTYpFe6YZf5yyvzxRJHLJ8U7HSeeR8q8xrknZ7dXyUUNZuZ4PUcutoZ7HnOIAqSqhaVirm1
0eaPOJUDELLvkd7y4gN3zLDYTcmpPs/GRYkShU1HfHrIiGJshAkEwvt9yj3EQ2tE6AA71ck9GLcT
iPttnDZqEXKNxzj3w7gwIwdJDZ7M9P4NLf0KhLpYA02p0ybPUIJqWdxhFYLN2n3PBDXDNbtxGqEL
CO8Acto41J0tXLLTBSrc78SsQ+KKmqOlq/EnndoUDBAMivXt904u3SGVOKalpNx3w0oNBt4x0S1q
dy5QovviQ8c2124OZvXN1TTfYRQamBTaTdH6w91HpMu9MtVhNdtjYRg6cDWvEarF7RZ7atEFa8nk
knU8o7wQoduV71rqcNr3I/PJeZ6KZQTeFZaxV73GuRsN1MGEuI4NPjir8kuNjtqJBV2Yc6xnc2pt
sifoeWFuU6chNFOtybNiBiDy7SfT46J18RUIg+PsYH4zaocViNP2/CKqJd75VrkuwenhfXfcnQ+W
4aSCVVkEeaq6AeWIXEfMUqLESVmn85MFQU93qw+AvFOZS/CU0Oeax/Dy4PosBfrcXYxsB1UxoLhg
stLt3eSDVWgutK6K61ZbJYHHyk7kfiOn+XAdmkWF/x7ghckekwJZIMMt3MlI11cp3I4UrqhC3YdL
9OewS/7BBiB3Ylt6bjryKGKPlz4CPIwY6qyml5q74zmmQrBjOXbhzbJnaUw3ZanQyIWZphKwPBzv
zcSi6EkNfKx3dlN+McBw0J1liEodvfixK4q3vDSYOh8EY6z79TgxRBfrD26PRwCLW13+/ySJKJYG
rd89gtkNIOijuBZRhOnrpKErylVt52nRWsqGt1dPHGBvfIjy1p8sv7A6tmPfnh9q2WOnDC1FJwS6
gSDk17306OQi0hRw5BnH8ucSqUi1v11bpxhE3JBZ1xU1Q6GRA2OXLtGeyDBxJG/PqFA82dD3lMvb
GRQESgYBjedgJ7vnxtMuFHxbWIunUMpmVKUO7JiZTGH4gMCh693sFLwjp8ZzzEDcBp6TRAEfBdzL
gJOp/5bp1L1VGaUdW7d2dbRtIDQlqITQ6/RARXKazY09jaClHs9ybu4w3d/+J52UQ1keeRmlbrCr
LZilHo10z7fRex78VIUNCZRAPP2oVF1OGZ1dICh5l/uz4Y6IIvF4Nx+V9GB8yIMhGB+oCz1kDejP
SgzSJtQ5E5ob2/fFjGMuC1SFZwC2+bXeiCcvc4ARnq22QA9UQtXPkCBb0UTJG4B4rklbFgHuTqtm
MARtF6uv9mNbmLkrAjxp4eMvOcz3vOH50dnHr5/GSlCDCp4VJHGydeiJHW/cDUD9tZ4/45V66rEu
RFdkfVQzQfUWFMKNNT0mIcscOkn7DCRt0hX8ifeRq5xGaaOaxUeysuEAFyntwupTpzoU1yIq4uWu
dK7RD4zUeOv0wZiHvvPwzVXdvnwl1CC+HWy8Yc2o7hqMpA5Y4uW2ZyFNWTIwiwNdL3bgTbcSK3wE
gyy5XiRPntALBRgz01EEUG0xfaxxL4T+JohxhhjMGsnf5lGoxmVB8lrEsTbBu1M2Gg5/tHwTV06K
bjcyeCi+fkPj4Lxri86XFSAIyNqy5l05dAE1jp4A9U9suTVvvdeljENTGRenEfe/iekgvNK6rSY9
MzqBCpY7d9M4UpEEfPcYwgsH08pRXReq6tfmTtMmuC2qcu9UKLEwmehqxqyd1bn6MW4da1T1D8UL
iRtGw1kD3iFHeXsB843A9SKAZ1VfRfT4GltewOc7+b1ZQZNUUtv+hPq11s63EqKNRGWGWEkqzrCI
63HWOGTh5vIZcdtuP3gOCyWc2PZz3YIoWRTiiqQvnS98CrA7WvskcRHHw5FFwEAIaZX6Nrf56MzF
DBkSUbOlGaRZNDFj8fqhl76JidpR5Ci5BeCMSfDQzq158l1vu49HBy+Ci1tM00yLENrU+Jd+u/il
7rnY7jbDlt9PE3WdoreKN5HSOxDyT9bLzNISw2AkD2KATL4gXYDNdNHBNhUIbYJ9JaeUQgZmEHmd
fmSN4KGtyKj1yPVSXPIltvGk/VdZvJ6lEpKNtyPrQMjouGi4C99fjwpYSwWIzSUQG4FV4KIGK0FS
/Q2h1Uz9jdtWB3T62kKiPomKauYl00bbIIh3FBMjI2LIJLK+ICw1MXC6yIdp8nNFqcjfwXjY3cSi
nua7qJ+hlbDf8+QCKP3Ii2g9w+D/nz8SDtipCZsEdZg8Y26PgQCiNoIwI/u9WHU4iBYMxP3epB4e
JNFexryYvXn5f7emJJtyryu2egK0XnFU+1N0/roK08HqqD2kXw5mrdq0D867XdT4quJPJ8T/Id4J
7yJhKYgiNiySqn9AMtlPSZ6bVOs3S6F6sPQ/ZsUsCwo95J3s2T4Cjl3GBM2YA4FEwLYLctpn1lGr
nDPr0xzYCWOo4Tq017zfDz6GtXh8eG6CcIyI2ckMla9VEzKOwSrmlP6XQALKudWYuDz48ZLRhJBW
eIg/KvWA5sQmhQ6Y0m+3WPC22cTTmsfT4pbuNpQkmaulLd8XnsWJFyIzi2by6CpOk2NG39LQIUZM
DK6UchYdHRz/yk+X4/TxrABHTN80NH2ot2R4a8TzOYzGyrHwDC+W9raw0ssKNDUChJoyxSygxQQO
dn86/CUelDcjHr0gRzCn9c2Tap8VLbcTt/JikAv0BSRB85NpXcieMsT6qXgxfjR+7bxef9gCFgXh
MSFKrXzs8fZ8Vch1T1oPbVJnWOkGHymvq71sFhp6jN1OUK8f0Q4lDd3P9elgSb6yoLxyupUzecCQ
10aoHXlSEeBbBTuosMoLfcZhTNYRZUDkiidy5G55yGqdK0KGrelELc9nb2cBSLQpT6P8ApmjAgdA
2bQD0EAm58ps2QEr7RzHeV35DrI9UYJmHoC0/85q303dW5twrBB7Zu6lqq4VQvVuJozbunI5Dv7s
rQiIChyh0bOpEcfEtrOo0WflcSVMOabq48GhYD9Z/q1bYhfhOVUNXrng+mCkRf0keqokLRyggJDc
iyH/Dxb3PO2ZQsAOnTKKBzAGuuPEcYZDL2rMdgSRgyHbRBFK+U1hrmI3OeiiWosI2/Dmr7w0rZBP
94MJbeKALAohulrQsPUiFZApMaH9++i7CQLYQniTNnZU3gvITeyQYgOkVZDeIJVopLJ9Ss7WM/mw
pLZ8O0bEtPvxcFkQinCeq3ugmllxvbvZ5b/NpVCx7SfsaX00lNcC25caMetjlJWb6gP0lNPJmnRA
QiyYQ79+XAprRKfQQNgRfPqI738g+MLZ2j1CV05ILseKqVka7z6JplhxrKpLFlT4+Cs6VbRvL7NF
u7MHy2Il7mmUk+b68ad8UxWtyBoiGpvKRiwAp628zK1QskIhG5L0WnJOP4HcJcRv4EmvA4GIUluh
bUx26McOVjDxZIXXI6iUMXQ0jjpbR5XHeywGwt2WJucowC0HeZtgCCakg7gdgKpUnpuyCrFm3/tr
R55D7DgNaiHatUcargZqK7JHv1OzKiQ/k/T90i91KgsHPI1AKzEh18GR6ypnKePgMpBcxs2uCsXz
sM5hwEaCcyOWes9IfOE6DN4B643P8luklBkRQGujlyUB9P1Nlu77AUtfxmMP0NneMGygyeGaZewG
uQHR3W61/cdlCWbH3SMbEwp1zdG9sCp0T/sRlY/zEO0XyPz1Jek7sKo7El5BBtJWv5mSKRwkO4TI
bmgDWf0qh6+4RfBS3YWAAeC3b31UFXp8QeXTwXD8pQuv5MsJlTM6VpIsb2CKnUYEMxv4cINbNh6/
EfaIpTHQGC3abBOsHtSSDh2lpxSkjT2TW0B7xSdljG3vPwCXwtkCBhXyGvz0Rz01wVSfukcx1fHK
WSCExiGJoCKUT3/Q9oByvavJ+Ct96lFgSEkeZi0WWs+BNEBqyhUcOap88zl/jWK/jwQp9w9xCaK6
k9P3/qzsYuaYEEFIZGM9LhLDd0bwhWvv94pLZc7XVYAwebVTkZhTEQGDq7/Qv7i0ogHw4TF9cUC0
UwOO4omZXpFrTKFOqBs4obb3JlDOUymPUCKOzWEvQpZybuBWh0Rhb9HEh+XrLRSJJ/dcq2K/+6e1
TBpdqjfqHZIttHiJnYm6cN+11oNLn3y/j9f/Wk5UeLQ7xUGxO+19TsEqBPZKfJFW5rFeHCNAKdHn
vPqkj5AUh4OvNeyWPAPtAjc1ar9zBj/Q6jskl/xiAqCzFhCDOZAVpQhEoQ8eYKZhIpCOEo0R7QSv
nlQCtct9bThmA5RgSpXc1BnkQdR9/e5GvrfDbgMq2sbmsmvPmXRasfXAb9Alde5ksih/kFK6j9D3
b8sussAiWqnlMiwcb9Gk89/1ZTX6ZfS2lA9dD+fplo508Sh6gimnsgVKMSbiBaiPDgnRV2LPoViQ
T7sFlNKKtRjzLFXSn3FR3H9vpRcfNuqmbd5XLNf8GFTJKUWeeRBcXa1dyIT6ad8o5Q4aQ8qkF0qB
gjJG2+dPRiL6IrkOOuI2oUXHe8DK8Ehn6wojkG1MafP/Xl66DbYTPBdbZi1VgbP5kcx24gj58OF8
+qKWb9c6cYB2J+Dpxl6brL+OPiIUGhMmVWTmb2Q11gy1c5QWf29Y+RQ0iKxZsA/t7dTBZpVZamUQ
5IEnFrfA/rxHxaY3fCPcI0Ph98WZvSzEbEIoTHpLa7B4moJwb/wmEjNE+i/6rSYBWJNDX9IHcur+
C6pGRlUIDNxo7JXPw9So3RImDSVbz3Aog3SKpLz7GWAWTFaaPqnKLQEDAksd8Hd9fVhTOdAeZRfm
etIGZE6BY4EIWIRfFwRpU4fLmnC/hzF9Ax0ea38EoptqOd5h5q1226K+xzKJazF+Fign6MnH9T8+
J/+fiVsiQd+Z7KphK7Kzx36K0A618V/Gy+M2ItbRz/UehMW5CGRq0r9fNpHzlP6t1aqEhBOXZzpE
+Io0wQ+PPCkuJj1lSbKZhJxlPJxw1uk/Sge5zPtFHOf/KTbTECBSHXd2QaYBD+e8vXi5931bdBuK
s2gVQp3Hn+vdlxPxURoYe2dqUsrUwqurWHTg0rK7B97trJrt0DtOO8FdA0al/aYJY2KsddDnUjcr
nlEPO4bDKfly4uRn0wCZXsXWAa7oZ3SePGo0a1I9TePk8Ib0glv5KkQKjZLxJfXFAr+nHkJ9pXRC
6GIRAfFvhWonTjDvzWtuLqg1JORRJ7/O7MvDEroyvFoN0hLXf3AxQjZTxKa6RH5mueqQDynTxKbr
GgaUaqgOT+5AdYHKQnjISFxaMGqMp/gHgsNnaqZr5dVwm3I/9hhYINxbUV2l/k4W0Eqt8haoNpZ0
E2ZtjiITtZWeeBwLgG0vCPY1oq3FaQFoaBjj3Ha4KdoA+ftAckqrxxP/LvCoHdVyYInmIacvVeK1
dnl11I2QAMDI80St/93oVoNdyvbYnA8nbg4/O42cLJobHlCMIGkIhtDxlj5ke0MKnNcqwXdIt7yY
HnLNHHv12sJGKzLF/+JnBtRZhCLoPBMzqWpsxBMEbkutQ6H26nYLN7TK9/Tu6focLBr1xQ0iqWwe
mss86yrdOsqw3R07vOU1qo8dCwUkaqbOHJIoK1P56s1Y/4fBZ8lTKPNtRbXxxDUmf7u146yQoy3a
sFTr3feB9GI0iPiYE/Qe+ZPu4TSkPVkL0RHKdz/E8FKh1Zh94Zbgmo4nn/zFFa0moYlTJ/P+VatH
ZXL9afV4zM1aRA1gIW69lyX0hRPXWx5T/20Ef3adtItCPeiZcEes+wVMiGeY2hy0JRakIjH3stT8
2LPjnzxJFGsms+zqqq2ihyscEeYAmxnzSZn/8YVUY4DizWXuYxO8ez0726cZwcEcQS9mpsLgWa0C
NW04Dm6U6eSkHGVgJJ/U48azwbQLL073o+VK/qkeXlRLQKu0yZlQmNHS1ZAaYmCdWIrFZT2mfXGJ
207LM0uWuTF/fXgl5yOkAvK3yGIln2MhNRPHGsDsXtPB8yD4/43eYG0Yh7WxJtCSbXtjI/O67ubU
RBzW/MSrr8MfYZn5JF7Ou7BAALP9rbP0kZGkUJeF5RGMsSR/UQlNZs49TK9E7VHX4z66UtlrXxOZ
wux2QFtNuyqv6IncMv7FViK/JX6NeD068JFPtoL9BAnV2pH+SanO8rSFDAx0qERJaeb3CmNURPqu
rifmLDcPjDWIlfWd+g9PMYj4X3TZ5v84X2QC19SDc+AdbUXxFj1Fbvg2XaxwM1xw3B9XXIhFiI0l
rsGBRVolbtqHrUFbh81ND7Vo6eOp5Et3rOsYNw7Nds1ZoryKISCSzpNDl2Y+SUeT5olxAnfcKi8V
x+NJFljLO3QvXK74260/42eh8qPR7h9/H7/erblyVKffEcZnQ/rtOnHMEkiNcb+ca3B5TfuvFNnk
h6nM44CwzOfStovfTv9ecVEEl3GdoGMpquf0oSKZ8/WbSjZYZSE8n/kYNU0+qCucjpAi013A3HkP
WOdD8wxsRUNAjwmNSQ67FkOCAOTBZu2NPu35A65LZxLpqCMF14GwDqyEzDz0neuXCaWRs8RGLMrn
F4mHUvg/xaXbsJ7wwMKbA5h3s4Ax44RxuoDrOXc2NVxcG4slCWJPxVxCZOrrtP8qw9Ko+XS8mRF7
ySbdpwgAKgV1ZHg4b71Z0YVCw1OCbGjqtQI1uEgkkcPlght4m8rGxCm5xbLBiyNKQ3hwsxmWY7+8
kVirRp99dfh086dFD+2FAKLhj8ItfNznDQACmoAx48tg++AJCVG9XhIsYHm1O3G5WblbU0/ys/cK
k5cNtoqFExz4XWVOnzkhnZqVwYi4/IFL3vWgOTSuylONDuSx0VtXXVkp7KI2bswgXGkBD0GIYeQC
/lG52YlJRxAHYaqUMqlNfbOqn3nNWMG5kvrgYpoDuLk0PfIebA3f48c9YQ0vmX42wRTy2kZiOrJA
PPq4rc3C3xTAgc/k4DDMWT11RlI8Hw9IjEoKy/hqUqggGfRizUTvV3+EFcjVADpJKEWk+uAjyMgz
b+/8SS9TqETVTfGtZ6NtX3BpFw1Su2ZAzB2OdlSscSW/zpxCnoQ8qDWI+Or2RYX7GCoPKQ4ZKMM/
Vf04WyoYOjBhQpoaxZkXjxa6VhY/WfoDiGfJ/aoVRkiOSrHCXy4EQvN8fZtsNaHnn1lCUd9lNHVo
Rtx/IX6UxXdReT5R8LOMd6BSlkWFb0xNflhGaaYQi+1jiN0l766geP1Dv7stDIaGilweVfRODXcW
7lXuNuK3l+ngz37iHQq4BiOspOWHYHFdlve+JX+KFKbLHJmPce3NbO2N6hkS/qYGg7X/zE/d4tip
+Q5UlXCLji1GY3rFad23OAmCGLMIsrDHSSS7f/FWWKzl5dtiaUE2MEhDBrlNQaKNnZIePsdKaMS3
s8R6wi7HP88QzxHygTIhVd+x1RkwIW5uapt2B5bB9ZSLvZJnyS/ueW10lB3d4SEOD9am/kAKhX/B
6o3bCliDN9rNJm/XlxkXBqB+28EWqC7Jn/IXo2xYUgsweIMxCHBaRdnFl9aYGAYmU2ydCKNx9nCn
Oj7lsGk+s/8ehAxRN+IqOADAX4t0Nc4IbmNfa/f+dXVy0/fKR00qNAVe7W7fbYkMeHnxn8Lr4pJC
yR9UEJB8V7/lIt5rrOnzeUCdBziW7otHIxdFzqSLlZvHQ2qVbj0m1mTe20h2N21WucVgDJlXT5+i
X9p2mAHZ99GhjyIcLsRU/fYFhEPYtlQmyDylHEX01maYbhpN86a4Z26Hj77LZ/MkgEVjXJbyJxlw
I0d7bONXHTfK0r/IRai19IIPBMMcOZV8ZlpG1F8pW79Mm26DhAPcbFBVVcAdnVADAEWe16LdhsWe
Ocer+f2+Gzu5ZJ6tiZEa+4jx01QILBM4HhhbD6sstyZolPqq11DIuxeEuNfe7b6QZDWmpXsC7cCP
8+L6Joxs4Tp5D4h7UPflZ/Vged3Nrcnen6UawJv7vT/vSFMFvbmRqiinu5L1v9Aq8NCiW3UzyQ/4
7c07svnQSgW0zO8sKXnQoIA6yzv27uUVZBfiWmlg/woE00te9G+CDBsdc5CK1bZMFZR4Ky2J7rLJ
UwRYTxbz0fHjClrywR0U+5fsHPKFMBO+7/b8Rd43ipdJYjNFQpB2wGTVegTEOCaNpTSPaLbBTk+X
pFNX9KXtolxgfmbAhLRxmYoQsY/bgk2xJjGUnkB8apxQOOZN+ULNzl6ZeTRCf+7yi45s2mjCkrp7
hdPA0lTHjDPnowAHKY6uMmXp9rp0/FhNlCqDCHpN2ZVZAXE3/7fChOcgKoAgkPI6Lc7BQ4eY0nJD
ogj3tKtaLDkMmcU6MOhmtaejWz+IXLEbnyTywp50pPR0nsGU1PGWlz5EvRxWk2juIZ7dKhW1Mava
ohstMx9bxNI67GUGI+o4Ti8RU754QKMHJgKkz5wsMu4QJwHEAhmCVsB/+dEdLOj6ejKBe4WMVn3y
tc5z0KaSGmDDnx6xJ5Pum9blk9kE2jt5l0VM8+8uFKahniNV3mnICqLL4a2aAXikAw4v0zaDe+Hw
n21ShhQTDKoh34TcenDpgfsw8nDHDIcMl2IonbNCktiV418uSAX3oTJXamObJFYTNWRmLnalHC9M
Bi00yc5acrWcbsgz2dhMPAqHhHlX6EQ10zUTF6oYaQ1DBlwPxnbPrtEufpWP1G9KlfHV/mTZ0fBR
q+JY+pu4WvVykfq8EOujW1xmZeYVUC+UwbiSeLzwMIqU7AZ0brxG2rggJ/x+UQm28oLspMlWHxsp
mo8w9EXwsIkBZGiYreKLGIaMNdRCwquhyC3kjVD4H7+ZPSJ0cigE7QnQHiPooHSqz7Pu9dJNJYo6
pVGr7Ym/oS3n8IXauny3C4TZlXwm8d8vyks1UcO5c5XxVeUwck+ucJvyT4lVJNAOwQdY/1Le2xyw
g/idxt1UaEjqIVYz13hPF7iDaJBKI64MH3tpMnp0BuYgztTj3kupG3n2n1dE9nI+OjTNfFZaJkj7
NdVpnzhosiipSmL830J2TlXBnHnwvX5ouahCWQrKjH74m4pZgg0LWOdasETvd4rWZ9M1hH84DQ5S
rKpaP3ibDhSVko+9xMev1ugM+TeOlaww0/y63DJbafPeRIG6hXk9jX+U3226PbbgDLK4rkGPwC9w
nWDtcaGNCeG2ClLetXDYj2hq74musvDhgQB/G32urqoA0Qxq0JSxgZqCNPm3Gfx2/jI+d7OTH2qU
jaRxuXeHjX1rOKShPiyLpAHqgxeGrV6AYMJH3gX9k1gl0zvJUfOW/84ITUYatlFKnoV9DT09XbW9
pV7fDZruNlvDBabHDerkHTlm7OCAaCFRDoZXS1oyfn6DvCahc4kPxZXyxn4eRyihiV24EryOFrGn
S4/8I4/BgplYLGZblRFEFSMxV9miD4Yho8q4cYbI9U2JJ6TTqRTfJPAlA/2X+QhH0MJcgx6hdhXr
NFupZOdCphZFIA3j8ZyIMtgsCMxzAw/SUVY5mTNrYParss7O3G8vGLoL/mE1MKydn9yw7mTANLnm
IswCjJfVPgaNbrlfPapKV12h6soe5phfziocD5g+7j1sBIMAfyTwsAIZ9P3Vzk/B15iwj3IVdD/d
xA6xtC2bBRh+DfcZRRyx200bKINrKEgfcXiFR+0w46J6QVix4h9WekhiK+NHPYk9ikm/FRPEBcfQ
m0Vv4LFU/jeKLx6dlFoXFzOgDOANoyC7N88pISQ/KOMR2fESrPe3CBTopJu0GBSk9WiJgWzQ7kyP
s9G1S3aghgM2Ba2xQDg0wTctmrkALuFn0MzeGhStZUjWJBQAgzL+vgHQ7fk05VOFhFOJO1nmhtG1
RLkfwpi/hA3dB56b5XH+r8Uht8MTzKm2yaG9arZdPpf5eh6UY3q8nHAbUoFYxAFhscZHfijGtZK+
goZybE/7/o637tMqeWW8tBjwJrLgpT/UrE1BTryDcdKi/UXLHo09qZ0K2x8DIVueJzrDpfBTzoXY
6LFXF+2RBjtArA0h8aODU+85qG9EXAeoxZ1x7BAvK9TSqfDhO/I320ivacggpG2Td75jp14eGO8q
yXwFgXU1aEdKq10c9rVmtNfLZXZeupuMxvsTtoGQXg4aMJvNiWrxL/qkIuWrvWEeKUoEDT2JFABD
0xUBZ5rZv7gst4lH/LBx5vnbZU4yTZ4wNnVwrvMNnSmKCNbeQXg9NcSCM1cbN5hbkUzo/srFA5Lu
ozX525Js2y9IDsBnoiAA5xlwQvBu/zC+4sFd0/chYSdEBCEl6SUbapyyx+fFmKDHjDRYuEf7TLut
S/ptLp93tmWwpNmxie7dJRuRffbv+istaOCe8JjMg2IhFR5PMHEi+rTfmcKTiLyq2goDtOSBkQZh
U1wEFXTlKG6OXMgKRkByyjaLOdvknmeVFddwVD3Ux+Cd1mFHYjn1g6bmyOnJkTDuPQLfxEbQOuAR
Dl9IsfOelne97A4lHHXAJ4KObnRwlwgh5MKXTc5J1O4IY2+3HqSRt9b6VuNoXfZDN3ThVJhd15cl
lLdl6AaHZUB+d6/KM/vB902/lW+9n0VAL2QshXPE8RDOjuG2tzvHpM+rgvclrWkArYe7oP7aUCwH
thKD7LC3N76Zx8nZjSnlB7dqnje2Ov6geugP/y5FwvghhSv6+/6F0fXKYx30tMRQgvtQPbwogOJ4
4f5lZ9L70O+sFk9ku5kLtzgEJhlla0uMRSaPDgoXgVhYuLzqVXmXUAsd7wGVN/UySO32lWk3S8en
KgCIpwyd43TlKWTpV35L/Y7VkG+jM/wRSllIxN9W0xeLE6zD4SjFCP+8XYQqgBqNGBYYyFecPlWe
5illVFR+FGrEI+zDZJO9GN6X6NhhqmFXQSjOVv0wv5anBe/h5reg3/rEzEFb6LLIeF9KFX/BxQIU
ZqJfOl8+rRqXFQwnyajF5KyVPt4p8Us4Pgk7EDYnkWF3UIg2UIp8fYgbFxACWHUT/nIqQzPP0mYK
NIM82C4cpXqZB8LgGJUwcIAi01+x8g+Epj3aTkOPJ5dcrTzTvHSD29jgTm8WFMVP83Xuq5FVe5dQ
OHVAx3TG/Pox52xgGUZA759fhYpE/P+f+jLRr/n3hZapIHxa9XuWlqBhfHa5ss2SL5mkEF0znB8j
zvJxgRug0Xt4q4DbDP//9n0hqMPnB7dEcetfaC8huHi9IxFDiFqjFYxr1I1u2DM//+D7fRM+pVSo
NMCtgpAw8sKjw/an2xCUPkLwSsMHhTjpenQsF8meQvlUJvCiVTgcVXPay7D7kq6dSxIARCBtJFt2
KLs0bQSukih2w3Aj0LDvGB+WnFNozc6J7OqYVX5rb4NnjUwgqg8gthP1A/9sSo+pLtVlhCf2HnOV
fw/hABVUkyOJ5zzlePesplG4xhwdAk2eiSJem0TFnnex8nY97Qv7otgd8XG13Ou5SV7MPvLi3C5p
XFXZCPCNjJjpqwdfn6OkdWabbceb8yxpVmrFvWo3c/uTE3TE6AyNnb3dF948xO6EFlXaq8EVkn6Q
tjKpszpfHRjN6g5VgHn5Dbw63B7d5ee2+IZEx6JovyCqN8LUBUxCrFJP8Tf9LBjSjwI0CnFtg+QI
bO9M6C0rh0k3SvrG67EpswxTdThkrnvgMFA8zoqMiL8yjraw9GGmwqV5AbvNoMlzyK2JRA5c0VIt
kIX/yTLh5msHOuSqd6WIAgAznwM9llMPujBPVGtlhttPqXWV9sENW/RAxELAps6C1KU2I4GTeQKO
GP2uq3Pb6xNh0GC0Gv7qmnbkW2bbocW9uffEAtk+pxkyTfPxTOs59ft0y1rsG9Oqyh04w311w8Il
QAxHdDU7xiswHA98ysyAW8f8612X45WOtVzgDO5nP8HISjxBNLJTFOX/xIwlnFt6roGrONJXdKPn
/xuymtt6mqI70+19WfQFfubPiv5Fv3bvAHRytEuOQ6lc9l/swd/2/67LReCO7/UjFQB53bAvFh3p
Ld0fwYIPDY9gaKyjqW8SJHa1n9KTtYiYDeNo1ua5sXFq/aFUg77tHA1ifns4jGARt5SGyntHs3WR
qG0M4+5xZ1eKc88RW5J1A2RxtOSXFPR/BF+iFRGKjhkg+JMVMoE3QzwiPw0iUjFCtI8HYyDdAjqY
EIjoAt9uOrfDwjcelBXvG8rK+znrBRl0OToGEiyvJb1Rfnci47GOfxjpngPLAexgHyE2yOPgpYIr
/8JbZ5j16IOZ4frQKuZvQ0pVLCYrd6L7sREBpSQsKwzbbtBX2pHC5qkLKgyS2KYoM9mrlsmTuad7
5GQe7sxWjzssk9Y+Cnii7k/rnNVD26PdpRqpi/MWdwj8jFDwmxcJgvFEDRRNLlWLYJ11sWtM0z0o
TnydW1sJjp9lSww5Ny6uq1SCJPewyOmH4VtR1JbbbpDvvGpFQuzyLS3/LZgrfPOF//HAYdVG2M5B
AuZ/+QgBKGEtn1Yv46dF9hy3o+ASbhTjRKwZlEO4lHNb1vipsBoyPRXTJHxuxHtUN/h7pvkcUVtA
MmKxZlM/sRflmGlBHpFfhiEOFpTn//fKVOD8p982NQTWbnfEl0pJ4c+AMXwuqPWGO8zcdH0+PKNM
SqdMMfaRIlbOnLnz4nX8NBIBIiQ7W9N2C9Lrj2r1WN1Fkbv3sYm6lw2inIgkYq8w8u13JdhiHpqI
m58118iE4QEQDhm7vMXyQId3ISl6Sbzeg1cvU26oq4C1EKlQJxXsRaERDlMXn0pD/6c87n+MQk6c
axyn8TMf2HFTkUMLxy/K8Cxgq5z1RZW1CNhKo9rSQqD/LpJYVjv3FAeSqqd6Un99D5mfbA0kZPA3
Imyz7IaVOudx1ffZz/tiQYktL6By9aTWVEDGMxdJh7UA4ejv/UPPPvsULJtEoVxnMZdFo79jQS94
iOb/+RGaxNnhb6CtLY/aVLr50FTaiXsweQFA8CYCc4CnkQYi0Db2xSB/03Gk591MucbbNFE8Fg7O
zl/1Mu4dt9VqbV9lHGCeC4B8SMHgNYxEr/y+o/yQltoP2P3OMqspbtuvhCM3/WwWK9QJ79/SU9+q
gwSp+gahuUQ4jY3Pp+TYMeh1mm8qo3ufIBAhipsCl0NmazieI/Lat/yyI1HhWttioKsHT07U8yTI
BE3axHPSPZEw5ePI3yYraAp35BKwO3aj7pkPVtGKnoPicFXgHKfJ8ytcS9bydW/WV2LRYnUMs0hN
FTvtGY/aJRFuBLv6iAcfRqkgb78cjZE6oQTJ+aAYeUvKAAwTKIwaUUAEf2LW9fAmgFsydqq4pSDt
J2rKVS6WIlj1bBdEaq8OJ+TAJPLkom/zG0eySq+3SlH68B1C0xVSoQmUbF+bOWJp3zFv05ghC3zt
Gw0F66c3YQuXAVUqo76Ox5TEwR4WZk9YIj6IBYyPSwPzTeEW/HaZI/rC+MK83113nbkrLb0RGCd9
4L/H7ARDCQ/DuMQJsS6hT1VafilbCmFXDNYT1R1aXAznFpSueIz1J7ZdImHIyPz0KCcnPqdIUiXr
Fzw4DTUGqG5k6lHwRxVGtMKS5d1xLWk5FwCs6bZJqajrQNdQ39oKlzdpYglJrAlXQsyA6HPz1wdA
ErtKiDmbxyJ2zS7YzGYOOb8BiPaiy6H0IwJ+L8+IDWHBQ9/UfS9XoHWYO2LlbVkHsPepVd35xl7a
c4f76ZLbvjTJpdBelaItqh30yncc5n7jgjigtfZUBj/Ou7JaSSkHF/3i8sBuzjH0lg7LFMnCjL18
4L49Hp4Zdroz/dh5cpDt6hLySeDxf+sBBuowjQlcXamm9VOcFVaHrfRIK2Dm60kAiNNRhKmbPJLh
Egk/+UoUfp1bY07a2lk51XVzf3npzR4+G01oj5E12Sq7kpk/kaeL4LnOStGofVM6O9agewJIN36o
+tgNYWwOVBec28AKbX+nw0B6+ZsU1k8YmJtfsx80NubQdO9tmZXBtEQyhnOIFUhEPgEkUlgwciHi
z/kBleWxRwTVf9vQtaWeVsLf45P0c12e2ZspHDNvyy06Ifo+/61ofAzcTHye8s1on25RfEaU8/pB
BgJR+PhU1vnutoWpBMse6q71nuHtmDiqgFTbpIDq4sZp4ce373CzNIb69MEc4Qq+Az8/rzCdvCu7
2CCdmWwt9CD5lylXzsNRFFbKHTNSxqCwxk3J27ZlH/3PQ2HXON4BBG9tcrq3uhga17IskqljAcpa
/Icn/VjeoKWZHwMeUBEs1XXRNZMhPhe6CXQD8QT1couF6dJEvtpv6A0kVei84gJXmxNOme3LkB5U
1q6dLBRTfW8Yfd5pWn5Zh8S6z+73q0rM3VgrrQA+Qi7K/JmguvH2GH+3YgoSEc1XZ1r5vUwssDuf
Gccx34ZgiAphmUpV5PIUM5gxaNW+uQCevGJqOBA/yVl1aXrA9shHvBsWRjC7GbpkxkTjFuoDaTXt
tvGNFjyMa48QDBTRj9WBCrtK9n5r0XWWD9mGWBbsW52g7gTXP/0164aLSFFgVdeSk+AwzgRsJcYP
CYg8rnWjnn5x8RfRethGEeKPL9sJ6FDfO+l+GpanfBrhdGqJ7ZmAn+WYo+5gAZylhuqGTOWKhTvl
UTOwTxEPszCu4LFUmIKIkCY2//N8qJXv5AgdWVh/VVvzdW6JkyTiqxjsQFfWV9O6atsupKa+DnWM
uBzn5rAhfBZg3sIRtcglvet/WX9ClS7YYhK4E1n7ZWP86ShWS+CTn2uqzRyxvEvJUjb4qAsnZeY2
J3NNhGRAVBtYk9rWO4bRnUkhSDEP1ymxvuX1TZkAw64try8SN/M902U57Co33LCW8aYxrYl4izew
9EEgZ5+0EbAyPNLH7nWwsK2LnmPYQ8U3sEV/SH8JveyADXgJSLSV9kECdMIpWg6sTWmCY7iUkPG0
rJ+UmVArP4JiZIETFGnAYLS2wePom/JNE08VIWKriGd5no/Np9JkRjZ8U5v7SqiARIofWI3TiOyz
6mngB2xWU7w7aVXLMV6aosWibmaB5KXZIuZhxaZoEVK/xthv3t2j9sBKlrg6mz6xmHr7xy0X7kcM
74cJ035crQuXivVJhtLEHoo+VPsB49SORtsqSmznSDX5oyNFXZeJ1R9SfTZY1w7YduiVvnJjaIyO
mxt4Q/dBWnuh/rQ3+FrThZDV10KRt4llBgvdFMpOBYPc55NJoVN4rQbZjVk/lsGM+dHmGs5gEP25
YWBolpwJ94KN9wkpmpq4J9Musq/j3gsdPoaVXcBUHSmSXxudjWbRz6ghbw3QVdRVBOi3xgcFChkF
ZlOXkw81u3pZd0EKd563/UjlOpGTEBHeOKHzaIGohKVEywqkQLCgxh13jsSKKp+48gqm12V+igmR
kdXl5n78aaRLCPVS3PSKjmJWYacz2W88aouwZuNF8tJ/aBXq+0O6VKQv5pSWDAbUXIcpXLknD9Vn
nnVatqemcGehsMiWkHSGbLwuLC+4998kLmZy1duUxEzYVdQWzBxFnSRm/hlmsBW6XjhHUoqPgMDu
8jTrPxd3BkFBaOzjEXzTBG7n3gYEB54oq9GVXszZtQRDEjeCdx4zXxLbxRO0+lRKZQxnJ/BLK/JA
gMvVoQTrE0lXWYIooi57ak1MOeBGTIbdFemUVPGDUA39F/OVUZLB0aycWqX9G1nixY2W9xiIE8Hf
4rF9DcHXcSahOG7vb20ftiiEzfPuZdAG4PeXxBT2nDAT0noOBnvJocnAj+Ij7gEVtBLIO6iG6Hnm
1HzvDtCgkrjdyPmwULDe7M4e+ZHNafZt3k7Jddfbl+rjAE5qYlKIRUG1inuPWMOngmp27a7lcH2f
wl8RkBnkDjIYyD+9DQQhHckVj5rBvPiBJFctTforqBtR71EvPt2L2EXrJBN5DNBG/vOeqk9X+BeC
ZZ7piJpXRtja7ILbjVxuc386CQeOXBULOf8YCIyOtwHD+1QYF3akIPdgqhBSnhhaMglqBh0PCKMT
90Y9M3hLtuT/6fF1i4wE5yfEyG1Qre+NUsl6/UPsZPOUwOMEg8zWupooqr+FZ4CeeWFPTWLW7N1I
/bBLjj491ZGwHuPuSbLrabz+l5r133OeVHK5i9HFDL1ZQ7lKbYIWZfPJe1UdOgzNz4od7+IBjsGy
J8KlfldeCEEY49jWJ1vouVEro/XDkvDO+z+eB2VkUO6tLdEs+fxtn5/K4OuVD/18PvYyftwQ/trx
MNhN+VDwto1rN44hhyDmwXX69rZ58Abl+29elHaHimyJQU3KkZ3KocSCfC7i0eWOCh3EHAAf3CUr
eHUj/pf7XwdMyYxOrvFTB/7Du4G3AO/T533MdFY/y9Z5k1SUPuftGW/tEEbJRRZZU3qiFuj65aN9
A11O2q1dNj5cs3qP31mYrkEb6feZmhMZNBz8nSECAlqIB9ah+pohRRtwQvauakDB7WxcZT13lRgm
d34jfMFyQC44nxP6XTm1DHkuSie2LzE8+rSA/389AP7Qu5Od+vfFIMI2Sg/LKFeQJ/mrZLiuqgQv
KcttK0Ah413HwOTQyE7Ta5ug9ehflqD0SHrbYrZyKSthnDzw+bzMa2si25AR69d6fFDU8xUu9uUP
VqHfGpJ4OSHXAgu6ta7fhH6+Av9Xwz7Jy8EiKwjblsUs0tEnJQvupKbZ8w7buB27n4nb6aENgKPu
1isEyKclg/b10e//1oEWU5z9Oy4LQAjAmWzJWIsm11msH5QW4A58FpMRb6WCKtMtkJKOVOu4WZTO
iiI8IGdnjoeHqijWw78YiZk18TRqrkqV3kkCJhodPio5uMDSXi+W1FvwU7QHiFkCF3UYxj9+4njX
nWhfBC2HtJK4Z0OER671EZRMLTFsC1KpozR7hn4yRW8WfeCdc/ZPOze8AizeWE8Ka2NbnIHfzx4m
4unQvYqhRPaXHw/5UiNhgKT1g1QkT8bRFs8w/D2yJLDNHD4u/bmcBYI/+WhaumpNsongpPUXkRus
o9kIGktbZQJ8McvYwBdQk/FUIaYwxCekJkp7BHAOp61wOvWtxKYRBbjRnQV/7xBYcs3EtsDuCiij
B+qHr69ImJm/y0krpLonl/ljXKNSDrWjqiSCBIZbCyVtV/zGZ9jYPu6hxbYt57jGZV2erxfinWYB
xdogRC6h62+aAaTgN0dYifQfr6MHLY7qpyTcIgTjYptEDGJj3FDwmk74kBy0G54BKC9eV7eWFsbG
VO0hCQA1NPV9V6LrPpmM3JP1Ub646OyB3cWlZxjsbsLAUjllj9tBo9XpM3SzXHFasEpzmx/O6uaI
f5/DSTBzjr0RoPiVkDbKN9jLjuG6ck3FEgSTqBzl/tDLIj5YLIHbeCZkZyQMFxkBJ3yT0ynzHvSj
K/qtR6MdfGeiIkoiPvVBtxs/SgFVoI6zQUMkPgZ5QgrhW0pWA0C4TQdbNpeBpUIioJkW+9qQHhzt
fJYwqGQFmRsllJpJY3wbjSFfw8ipK5OjLkiMRrBejbFd9QhOOEUZigW2jjB2sZx8M+fW1MALENCH
ymjYjNU/c6s3vZhm02op6URTrMCufagiaH5ZmaqbWzqf7urqIy91R9cyBS8TpNe/VCee6epp872n
GJCIv5oLSle+zgFxdHyJhgoCSVsD2bYYC7A2+ikZ3iI+5D4ExSRsrZKaYEcQfYaq9ooU9TkGOZZT
9QK/g0okGbn3Nns1SSwj2qwNe1S+vAUajZNtjqOaV1h95wN/RGfl2pjZR1Jf5f1kiFI5mGlGjIRn
j53eYWdmx3mUyj6F+T49Jh5pnWdEbDj71tZ0pL18loGL3kjKfoHNc4ZuxWa52mF5POFF4Clyc4uE
plZLVRWm5SOXQqyAE3UUGIl9Sh3VlUsRFVlTDP/WVfHKtO9w2nMowP0zSaKBvmKByni76cc0RUHF
RljC8fKlK1m6Cch2s5nRgrTNaMToPa+ksO2lScRrkrahWMDCjgJU+9y5ONJa9q5kSu2dL9RK2dJR
dCTTN7WRe8rRIs0G1H8JiXZX6tYY6rj7+zgOgySNZlGfF8Wd9uumkiFr7vzV2yPC19gtkHOxd5kI
tPfBpZjxnKxqyIS20I05ruA0X03TdTGIU95Les4TYDJGmjWzECRF6ebp0zAIbZ2RNoVkWaR5tyyG
6yqlpBCHqHKMa/pBKG/aHbuHlKZTwraRvYzkSdEROHrgpqsVCBRegoBABxZTVIERlyFeyDZ35oFU
4/NeNG79hU7t+xILr2dn4TFCc/zZSEybeNXAoojOrHkWBnACEu7mNaqW6tvEZOD83UiE74LWjrwx
zvtt1O/GYDrbtwPm9A16cWhQHQaCJfr8lojD+RX5UZk1K2LVYL3tpRSWnrRlLF1UaTirhDHvzGWp
cvuN+jN2DSlfIFr1nr0CrGviQ4Qu0+0oKLqpDt6jll4L92HgNWE9AruOQVqFvtFb0aYjk/CRMY7t
Ae0vhor/xLNMEhzbo1oicl82hdMfzMWiaIja9cnwhGRLYgdkC3XmE8G5O/S6LszLDOWKroM25L/O
QIKaaTK48qBBlM9qVrcX2UONkmRgdwv3C3WmDihywgDBbjTlAJYCSebOz6dOBBK0Yxbx1xPwVHHM
HC7hLA13hlrQjbDRXVuhK2cv0QsgoK82k5R38LhPUavnCI4ZSW2cnkQT1UENMGD1CKHZrGNcOIvt
fw+vP3ULs08DG4b+9oHVNu5Tv25Yae+RHtEJ9R87QAoJzhLOh089vyHDet6rnJwKNKoGtevf8gkY
lZLhXgARTtNFGKAYwYS1oOGeikVAZC4eLYCiaVspvxOGDaeG0pv5tFdxwFkPG9N3XMZWwpzPVscw
Y+yWVoVUdn0Y80FYdjp8TXNWwkUVqDU98HIYm9iwn1kEf7u0dVoQhOVe2XiSY8BkMicc1GQXSz/h
ymd6uCNeHt50Ewhsw0bUkD8Aci88azcWkILjvXVxD5TlTFhkn5MptF5G4M7SDP+sshl0O9vxjO3V
edG9jknTa//iF7tcpO5AuP060GJqQhPKmMSB4zweDfRPr2KiB5dzKJrv3R42gTEWOECmIt/CvA0C
6yVZ1g1IAOEOe7tu4fBhCcn7ErSD30Z1taRjbSvQT20Axo/5QvniLBLNg1PfmdGiMRAB4f90aqkL
pTRIaatj8R/ggVSBpm6v57buydlZPngQkbrJJU9qqMiGZlpDlYnoor6mP0EDnJ2PLQHSolXJcuLi
9aCyWzINpdD/dcpT0OKOwdhkzk+iUFxJkl5DGtmrJX3k+wo+YlTwNk9hXIbIgwf1Pad5yLiewqgW
Tu2N6cUOTJs7ngZhVK5LeUTf17mIOIp6J3W0KA77Wc75I5YmrfAX00h0CeiT+0Ht4e4swvWfUa04
3SeQWrTAh1vrytwDgyDwkXFUxd56C4WwFrZKSfLae8d5IykEHQNjZB7mVTd4aNOwj4dU8+AwxbCE
QN7flZkitvwMhn6cNFvqPqLAePq0+k4H6GyPSo4COoLhLfQLG3pWgILTEr3mX/CY0IingnKKGpxZ
m1/6FuFWwmpDrNipkQYf5rHtrZxD+ACCOq9ne1qJkivKvC5lphDfzfJeX2I0+CYzSClBh6kChMxf
guGNP7F+OhfOCjW8aH52hwILDrWyOzdNmGckOCgWkgyqK49Nr7cVhazt1aaf1z2iGU9oFgqxdsSY
DAfyS49BJAL0wcbNpSooHHw/h8+LRJkS7N0YvYmVE90OlKtKfXZsuPifegjeftGtai2GuUSbovq4
u/wkKX9uZQigJ84VoewgBH4TdnB5oQt/sLg9Vkh4W+NmycRmxU8ETaFQ4fYnuNYVIhiJF0mUvHRj
jnnDvCJr0dbZ9udf5tV154xq6nKN6B1vgMQBeSbPrNpPyRDA9zMobsw6tZP0rgart6BemVFufDy6
8RZw+sY1sBmU4gf44u2LoAOp3FFcnsiw5SL7VX/iLRdn8pV2QXguGF0gf/aXyLq0nSSgpxOt2r6Z
tCySt5m5ogz1SZMsuXn3KCS6XlgSRKdQMFSlxNrRn+ztIN0qNoR2tPQ/waepCgTpxuFbAeIC1duX
yT1Z3qHkH/xvVcMJTn3+hI2IwCGu2haCi1h7gArbVhCM7RsvlXHZWVqGuesnlfrEZUQby5Rt86gK
Wj9Q1Swmy1L+VgBbzJ528NqqaxusvhKMHTO6LM64PNTQy4ubmaS3HqmtQ/VkTy9v8kYzfDeMnBkk
kyZfLTcrrMY5xvioLk2DRsLnPI+3sY+D0g3rBAkEpPNWWUy33UGivbtBsWrr+t4g1KxgWxbgG+8l
CsY1ACqZ1RgZkzUtUA5rlCLAn8Y3X5vZ9v1HAznsKWd5bgdWY24gNJ0zNhq8aw1kPThz5xNJQKb5
FWTi2AfWzxekBg8F2RdfHN77HJP4JFPB4WRagFEdwHYpY4wYnNhJTMHUWrGDwP7Yb3XJPqabppNB
rpoukXSokcB2sceBbrKau1L3OT4jyLMI0axTMqBd1//gjBcjenTt2zQOdtGlW8GUJ64BZzjH/Lmj
XYSTcvWK/mA+jYaZWM2AhsFmhv7t5BChKbj+v1OvL/PE09OiRAMmgay7P1LqTAYX2lyxyMh/bE0D
c6OXU6qPaM8WpThCgEZc7NVjEYh1V+vPJoO0nHjDdtLPjZAFcwudmbsnxvKcXWL+dNlXKghhZfts
x504TdZf2BGgqEnMgbdpKoO3qYnVZU++HvN62PjQigTcgnzq0eeNXa03O5YgXhCGna+uKvLVrDLe
h8aCR9xyQ88avCvP96NrCyLNGIlxlQF0UL0IoOcPnKAAouCMMrbIacCg/4bPfF7itDNaVp8mhhBc
lSqtu0QyyNsWxEUaGNBaVWlR2tF+l3TgmkMbDlTuJAvffZGXkTUTqjm3hYfEZrCh8StZEjFhFX1Q
z4a5oy6IRHUviFQoJAUq4/oQF5dGs9DjCILHVb+Q7AfcbuNeGLy0nFef3XZWEklJLdJclyKsAwg/
smNtdc0JYzLZq33IJSociPRssTSXfzCMEAffGZDX+MQTTxodyy5gqKB7RM8R/W8xTEEdYCDf8+XL
XRkgRkCzXd2gjyv1m67DCOM1yUUdI0q+F2sPRN843JlqZf45SHA7CdpC8zxR1VpWbNteUWJD6fEd
51QIV8NMCrqqKGXeyiCO44EG+yM9jp1ueUl84JdPaHB2TqeLWRkrB/HNaXE9cRffKAJCeKkd3RR1
TSLKvNMNkSmn007zGom9NRm3Z57jJvztfirasx7dhfWuu1tNRS0yGzZX0hm/QVPHfB1K33kX7Xxk
VntKwzzWmT5KIgrn+iBuvS2EYqOMhyIfIe1df20xxj/58L1Hygou8hihX/8OLCnAwqp34iP0bRvn
Uf098BNXj1362P5zi28NxjdadBNbuy5L7UBAxyfl0/DlEgUSVUydy1hCnEYRbNEUR+WwoaxUMYSL
LLofL9GQLRakz+YNourswvEwdzgNaV3IjoYRLWEwfie2r+W65CAeOLGcRequ38GxHH4XYtTNoXqb
CZ9qm9A5MsjXaD5NQgFgJ1qNFHZoFXQAMOpPFozEiKO3A0Fp2I+qiFppcTDb3yd1TByn8YHhcl0X
j76Cx6x6Q96p1NClcdSFIBe4AaA2YFviu5SRnEe4hQ+jSuYSsBx+DOoedUi4Gy+TAerid/ISnSkw
WGM3eVnPHCr+Z3kWZHTmHGujNTOqX1CaStHAvJ7Qg2rfcnxCIusTVrTlSxXks9SYOLxDhr6ikHdB
fgjkxnGA66hzlSh4UNNTkp4ZA+rnRJknOFKhhjE9Nb4WZ6AcmKtNIe8sz/ZlmG/GcRyPxZuB8Q5I
4ebA4XupZ8yx81AlO4Q6YFz0otxa87G0Fy4APCRL+VE755zEa9aSCpDVCsOsaps/AuyNeJnlSxGe
woGGO9ZP2iNzOxDbsbrXijfosFIT8RuBhfc1x9Oyqhp6BK564VkAt8NZB5nDi0SwDzEHtRjyNi4X
tavvzMTLiEGys12b8CcAUqqlx1r+4HrYNa/FdP4XIJ0/wmP5ssM5siCGmnSbKe3QlQEIf/SOG6a7
MXWLGxjuKWxeQ7EmTJUBcHaqHxK8QEdMGHxwXoV9QRYUSNZmBj0ygtHhEf/zxNB1VOCQAfvWI1OZ
yUA1ftwjgHP96t1cmrDFNAYAil1QpIvXIQQLzT1sZ+A+MYghlzaK+8Xt/WSpBnHzOosX3AjXrzm2
GmZI0LSD7VsyXJuS5dtdeIBClIPtVNWVCp+DblOG36Bo11eU8puGYZeYhKP4JLuYfgvOBG6IDjLn
ijhRqI3+FnkZbigWrRZga2OgoJvUKSqJdQ1VDRcxsqCDnj77i7qv3e1mMdSxZZ4TVhHNDY8v9jMw
QCHKjmOf2s5t0nKEoAolUxp/CVXb+VwQ6IuSeS9CoY3Px/y/05zVCEeqMXHLtvvSgriGZDPPPRZc
/7SfxIcUBVj2mIBGN0wf2LKtU1GH1FRn3i66CDdneCT8FjBaMB8jTM6PHwa8B8hB64IUam5aqa6Q
gk+NWG0eoDEZ0FIQTRqMzPr2lTpHRdd42hJUrnwatGC2mxKpY8xjXpF47P6k7r0ilpgi8vPp1LOF
lztgltRajOriYwjePxm8P/N/oipx3z070kjFUlmXqXrgQZBcF9F5z1azwvw86roLdmqV5fGEJSJF
NkvOAAtOCdgPr0EmS2E6Ikz3WS1xT/ZEi+JHKfD23U+GkrSnrBVoygzHpEFzf7b3MTuK8ELmuy4D
nuWe8PcW0dT6apPChUWRkhmDzRmnWvTJ3jrJEJpDBSq21pKdVMEengaN/4UyyZePB1fphD+EJ+hE
+7GDf/C514/T95wSuy+EK2Vww5Cr16lcD5/3k0477FGIqM+kEUPSVBr6RRUQawUhKlVYa+oR+hOt
6VjOlttoj9JR82bCBkDh53LNkhhNnAxHWIWSJRozfkJLrcEPkzJuhcrBSgMoMu1c+XqGjOM2VQoT
CRRvdzlo0Z5ezVroZvfe2Sr5eEDR+bw9ESCFevpy2qRtnpcbpp2t2Jz7A63eUkO4MbU/EGoyEqkj
2yQ2uZfygmZuLz5veNWE4cQBQDYw8ppPKj0w/9WFO5AWs4+veEnP25s9lE3Vw0hVa80eTH6HoUCj
Pgn9SBySF9poqlGoaB179wTR7h09CT6cNh65JUTHLOeByEp+PJFWSkzuUjAbhNpkrBHYk7g7Nm+f
tTvm8/u88gq+ocpOEuRU/KakcibHWEWX2g7BOfXIVUMNAI2HMrQUgPeTTDnOFYmlJcaZkK4642tC
sKP3h86Cq9aaebzZ2JHc63JM8kH0cGC3IBYnn/8/qmG2iEEOynVQ2yEXrM0qkQogbB9AiLoPEStR
xJFIFwSub6p1zzyDIW60PgDPbcPGyxFSNr7TNWz45szgBL1WJfDbOi2YZ26/KWDLVpFm+vDGiDu4
9tJ6oWK5RwVpGdLKVfxvAgGzFSQtLBd4PC5mN4FN/j7NudVUefenq2apQMk1lqQpGdvj1HioiFDs
HhcgF1N6CYmfiYi7m4s1fBRzeCUsqRUha06sKr2g8v0K/iMO0arZHnJ79JCSyPUCqZ5LZt8OkvDJ
yrO8GvZ211NYDQG7nWvAFaXnBbL4xEJjUVBdxHsJelb9SBqGwxAVStWa882KnvfO/miInmr3L7TG
ZDeEgBNG5ggQ9qUW8z9TVBILUxv4vsbky91B5uzBEgLFDXWQqL662v6wp9+M/pqYi9mMe/La1YFv
x3KS2YX3jDRI9vFU2QcvNkz7M8Hp3FLXZAA3MnBesW5VsA5pFOTGZyP7knhquj37wZTXCCruRwKm
zevCIHi/TSt7nSQS1XdhA4rX1cfWiXMDmWZefojU5m/bPIxT059PXED4AE7zr5RV8U0lvIoNxoLs
rIer0SjFv+cF5Yguq2xvo+xys/gO2GGtC2wHCu4PlgueS+7fsPRFhxK6uwN1WlQB7E8R5NQG1DnB
9HYw3/CcVY2DpZhg3ccN/AAuNr0FfFS0QPvHz9X2jEJ1yxUE75Sa/hOV/dyHOmEdi7GK5Mb+6Hij
ttBnqOuhTzbBOq64dAW6cgT7U1y9w182CY+aM20bkwGTz1nruTh5B1V5Xt3qZ7cHBTDfRX3GCMOu
J+l7ZjCzrf96zoG/by8II7MtHSDBrKPe8IS8X4oVjl2KfOFbtxwu5peatNqHs4/ZNVD9R3OrPUbZ
QBrNqAycuTlTEe0pgH5CHtzNDeqSQfxhE0pc0QaZhfpz/lkdNiOoCUAle0EWQxxiE6ZU8/z3yfDq
IEHiv/Am9IL9RS0hxrRv5RXhMUavDhA3uo0BGLXRU766CGMEEwfNi1rS9ICisFiyUqrpV8IekNcJ
vJ2afJOKl9pE1Q6yStxoMcbsXwM8YepIkUZCHKiz0NkQss90XVdp8aQp/z6ry6iKvXaD5aQNar++
k//EsMJRN4x9ZmIRfN/6/sx7PXqw0UUKF3L5YFtpzSbRvBjf4qKgPlfpPDJoWgAh48LNv5bRlIaC
G5QfIn1NRRHcxtKZP6ygdU74CWtpexE0P2/8eU7pmXUTOOiqM7yAAL4soC6d6S83CfZU2QjuOkEt
rV0xA7tleljg4u8jN6Qq0U6WE0I7I0BnPzJ9rVFCHRMlF8FM3CxHnMFcblnYOlH5eZL+IpxHecgn
AcQkysz5eTjABaSv7w65QAQBY6BslkCG6Lo2Qz4Haqxe7OMJlFDCEhC8bdqmFZosNWJiFHxNQe07
LHSeiL2e+MYN4PEP7pYZRp0O9WntS0XHFaJHH4zeGK89gWnZjFzCqaKacJLklt2NDw6bGezY79ZV
upo/p3xRD3phvCYAH8WqDgpmNquGAfN1zw1MMY4T7d8QXcPsntAHJP7fy+hdO2XSNd5RnjJLF9P9
6cP5qFnjpcdleIGeJXyUWT2zY18j/vrFBs+GjtaIU3XeZgi6k+Ea4KQp744IFb0Fo+0PrDMkkI+v
v1B6NV5iWiUqh013oZepX0xIDnG/j+hqYLAr4qdWdZD3ZWltT8lBRMi7aGoVRxFt49Qs7vc+S1zv
lnKwZkXOLKZOg04kINxvhT5tNkNEk2qjp+8zNbQBKv1FipvwQMfFveG0xBZDGpVHx0ocJsjNpqvK
REgDNVMYJLWRTIRTRWdur6vRmWmOy7ckOLHjl/vFN4uFnyYgNqPIRTRS8ZrbNFuUCPHbf6RDm14h
w9cDDxByOOU5/k5rjvtSdLn18gK4v0CTMbz2pKEPju7h1RnUbeFKmZJFyC9iR1Aopz0dx8mUCbz1
Kws3ufmJI6stxmGUujRayabZ1WVCpV8D+sx58jv6s2MVDenKJ/CEGjFKZCoOkmoTIvryWVxbx3GC
iFV3bltvDCUjd0ppW1HZHnwjHdiHIblk9QxJSWnYjtMMxrtd89Jy9573aIFMI7OGVo1CVEp/4v9J
58lXYSPWGdTr8c9VkJajnGDuXrAo2KTecvYGcIoCip+8LdKO8rASPtFDbSvasaaPy8mPtgx3wnDe
3lfleVrmqo4klHBxIbC+I0796ks4H7uenb233KibOoTPj5cSxtuM5wmbd8yIl6IEwprmqKBCjiW/
RqKuAsDxK8a+kaDp2r5MYoYdt8rDp272CJjQnkEOUDEE6TmmT5IThJwH21+6HXe6/4IlHqNZX45Q
BH6hnJClm/nl6a8QxT0U+0XkpBjnZTJGbqFG3kO8E1kxRlOj70GOecT6V+L0E0EvTzSqsMmpGnX8
CYCuqyXfJJN/JZ7zRkae+tmoC76169/PPMZlmcxnMA/l2BypiUSpdjzihdXwotG3bfsGu8FxA4pp
JOf57IKX6nnhRDYv/ZPm3VDKgREb6sZkrEQ32TyONK/Ch0P3zHbS2c4jOx1tIDxXxqytoDGlQWFu
Bq2YZVNl1YrDf5+EcyZH8gdJ5KCQLo9kBMLljuuwcmbFSmUZBdbhl+Z9y89De0fPqn/Pr+CHCgwq
VwqLtLDpXWUv/Idfit111dgxC0YEeChu6vMyHirxf1iBbVETkz5ntU4E+bnWEWMn1qy6Elq3+7qs
7idOiTayL3XPAP/xCsQDYr0HdjLlzZm8CVweqKY5wp/AKjxgiVIUv3yrIprp3ziyF6XsAQHEtjl8
RGqiGqBDtC9pryZWCyuCX/MNe5zUrcK9DyGnyO73PXMklNJyPLQ8v7hrOvqWYsM7M2jsOh7Rg4Zg
Bg8sBCYIKjqPJoI0EsXRLzqWcVt52aGJbXxUvF39BGA9lfoio3Q44AVX1IfKa2ptTAkKUucB0RSi
hL45LSwrp8XRFSj/nbZAF22cq/dd+YrzQh3KfE2bZ68ee+1G+wMeXp7TaIhTrQNNgsbMTFzOdPfj
4S1jxXgx1Y8uk9820wH3fAgb+VHZzBGq3mzKz07yQLsRk/KvYU6n75CNSNu+IChCmRYKzEPJAYN5
JkfMCf1VoSjhf3FruQIcMzwc/8/Qw7rW+Efh2QpzfC/Mo6oRhP8qLsGQ3FDw50MH+whmEDygxKhe
QfsqOYMJIiHh+tiPwPILq69UviA4po3xeOrWLzGVIA3EY2NQ9uQ9BCa1FabZIKF2h+djd3mWqwfH
dbxeVvXCLmgqFsugvcjk0t3s0zx/y6/oRFX2mYnFY0ohqaAa4eDm+pJ5MyXFdc3OKkhThg7s1+ki
V/8JtZZQufMbwRqQixGhgCRWpqC+/ryORjVGsXmIA3oySdM1y4dCXMbpbwwL0VS+7muRQf4QZqoZ
mdBDHnofP1Eaxt1JTr6Zst2H1JHaTf5smyI8jj33E7vep5la3HysY1eVhq/3t0G716invVYW34Ar
hlHMgU2e+UwhBFjaAtvU7C0T7AlRqk4O+Fy7Ksi3g8D9VW0XcEw1iFYB80sszc7v9ZJ7JJ/86gRF
d+BzYZJ19Hf3souclWLT7lLHS5POpZqB9GVT0c5l3dKJC1x5tF9K657LXbP0uNmBzQ+v++TmKKFh
NOyCN7Qv5lTtX9AVET5mmrgm4B+4Hfcf04PQE1QiWhz3jbJkzyuAc9RmpSDu0gTfmx9fvBnE0Kpe
UOMBceWlVsCtLpfrqxhnWnOdH2Hk+7LVPYe0lMyp7tPaHHxTeRf/k0qyuYQzdL1p/gTzjiFi+e3Y
7dFtwMktXa9coGqPIZdCjpGt+56GKRY1Mp9JlLsl+GSYdF+RmMLisOHW+f7VSrCH+BiC9EiPf+cu
umvl2ida6M725o0ILkwVWC+N+k7YFSvj6zE3IVkOTSoJ1Z+Mi49BocV/JAQTiHnc6ZN+Udi7IJnj
5FaPSRc9vUhf5xfwpSB9PH/3GN9Q4q6YKMkAOlzoqcw8fl6qTZSuPEoSOM8xG2T247CJ1RZ++KvG
fF8RsQ2UC7KHjMLvNn0GT9seSapn3Kvt2SazYC8lCF9ta+InNsNssUqrDr3u8Gz3kESCKSzfn1dO
1fsu4WJUVHVsd94HpKL871TmqxqTx6jSFjf/cd8t7IRzyMXXvxTN8HstsOi8m8GOvkUukzAjun6F
NAjgvneJGPR+MBAPV23jiauPmSKFmxLRpLgXrWPi8sQHOW1VzOBzKJlGbl980NTIc9VsNgOdnxCd
I7HMCMxgyDXNkwTUdTrzwu/ESVBOpcTypBoiQxk6IvF00xH8OCbRJKiPpH77w10yW1c+IwJmgSdZ
ffTs+eZFc423tLVoTiY0cXAl7+7OTSKD2AnXkZhg1xwFDI+myUURV668iiphP0hP3bclZXTXVhUX
KxbpOZDzOWq5T73toJuOv14Zl2ijGx7cKEcrTmJdKFDXNkgk+k/RPepM3KYGsrRMgDpkhvtFKfDC
jkeL70GxO5a3br4Y6swn0LHIPS4PqdPnkpTsv6MWoXJoJJ3fthKptkbeWX5QDQKWydhZGfpm4tYJ
oF/1Ma2QYocGwTUGB61AuzZjv4qLB3N8/h2nj5P6ggHfXMFQpGP1r6KjlMJz3PPo8vDjUnG4dFr1
rCe/HKtS/ZxJTbIPMeWVxfe7Ta5kSBIAxHm3dJXm7yPqp0EMUy16U/N6xCK9LpuG1+Qjfv3zy1OS
Y+E9qbCRKoB6Wd9FarhStkIhJ5JXP60NHj6SpbRJNvNhzT2XB3BJ5pFKnVVknSSlMvxYG2ZbeKgV
JsJreBzxDLVEb81v7LPbelPlKF6M62RyCT3oOgUH0Dc/xkuiqVM4YwbQIZQddLba8w4UJnx9mjz9
7qHcJKYdER4MDVSqRMBUuRqaa7gGsfBRpjqbo+/LoXtVMYnkIkcjBsPyPmzQMswovPSrg66Nr1Wp
9N8xBCEWyVjZX5EzwsmiGTqV9DPIagNMSVwiMMIi/L1GcUbvnqa5+y+dUUXcEgOHtzvBbSsUnK1O
AiJZ8VvECLv2OvMaIYCPEEGCG8oajZ1L0fuOIPxQBomuUJ5SGzpAS5VSFUObUhSAaT/0rDCtfQGc
3mtD/1ahjCEumSY9JgFHdcuNk/2IwHxKCnFfoOaqW3CpCh0Dc6eHKslMxdvhOczdGVKDVlDCfrOp
Gek/zrWyi+30BMiLuBMoPg+iPhin5uVxYQCzLhFDH9qQv2MD4uscPpo/eUl9+Q92pBMjN7FtR+BG
usjOSu9PaO3mt6A6N2sPVbOsFDGEzikH40DutDELQYHQ13vSAdeDOSuK9ZThjXkku6SQ9thHbk5K
5XxQl5aipqfw8g/tni1Obe2r2OxUtwdpdlY8kBDh6euDVY2qLO33EkskYXauEvpIZLgODqsK5Jut
S3hhIZR2/v1YxLh+gzHF1Ffr99/LgYYVJw/azI91S8drXytBKdHx9uUGA0/ptk1zj7ygg6KI9oXG
WjMDqdEskXr/x5yoDf2vsf7TilwKO7neap8crRm3cQkhRjr6phM62isTaB11Kq5YrV/5+zI0vPp2
lWs4fy7d4rO3V7CTfadRl2Kt0dxPyxsz6Wx+dVMWhe2yX7ZUZITqQsrdJcqcHvPvzxbs/3/x0o/a
vo0QxtjW2M4HBpops+f0ShiK6A9vyIp9tBlA5+CbPsOISgyvAI6OBvL5VrPnKBFtwkOLzkqDEoTM
X4s95Z4UrL+UG7Aj/LyvbT/sYfxPiaToMwv/1W5ZkdEz/8zppGdGKns9X8GPtT3Fg1XqSIihTsnX
5lOn/A96BA3Q9ZWu1Xhv3cTdazWTQxC4zSXlRrwvGE79TS+FbHrS9sCJOlCRLjrx7gXrnPZtggHT
kei9zA/pSMeISrxvSALCpd4PklPJVdPA5JnyZfTIcXA1jPVquiENQgssitGNNJ4GX9mDrToRDUx5
5LWLBNnstTfIY2DNcU/b3jdOL4PIfmknuMyLBxOKEDtHWf5yEq72Nd3CSM0SxQ/vfuoaRRL2uXZW
2YqCp8FUENda0/A35qJPFueScYmYAfK/32NFZdVko+arH8E11e2RPAiXoceUyF/FiTNBstG87EYh
3f/+41+dXIKIVnV7+ENw0De/R9v9tn3Ot9f0O852KHIX9te38FIJCeMpYadexv8uYgyh6yt7+36j
T4tTO05p5EVSvzoDMf9TfHfFKTfm8x45ojcXX0eKEYCt+De39w5sTCVXvrhcOcXWo+O0GljTR+1x
IRlonSLsGRlX2YGLbxdmUAJ40Yu5D7A7xhhJD3nQSBQ61Q/GmlGKwqZPkq8HIzo5lckTgRVgkty5
3GwKOdbjpNNEvUMb6CY2jWQF5F4fT/zR06jnBG2IZx2HksTpeBIm/tGySArISXMqNWpGIAr6coq6
JMqmMrbrDoe8m2mra0QPPuFdPpektewda+GvpC4U3ApWNMnZoAVG4X4stygWgoT8/TYCgLOTkGpI
9MQYLJ9WEEKYbgexnK2vCY0jTcMYuFgwRdFN5zc8qo1idcwQy/8tTpgPpLNbEOsRnu+uAe84Gra/
SOgz4Izv1Bm5ScoCtJAAbQMtL2UQlzMd4lz92BzJx+g1IaAhwodEU1t/ZeMS7TqnajdWCevJQz5u
fCeeagsPReiEKwI7GL0FzJF2J+y7M34HMofBRTrw90hnx+85XJQVX2crUmKCS0uksWlCtTtMty9r
BZCuCFB6MpB/msodOnUsrJJmz0GXO3ziauSGnz0e++6fYcvqsFzGJxMmcIptifZhYbyhfV7INLQ5
xTMbmGayK0R3W9nyFlyfKdq6OeV75HuoU6C3ujS2ApMobAs+1+hVVzUDw1Lq5nB50Cq5Knp4i/Jf
9cL5ZHpgLbjCo0ZWuaW1tAJnlAA7PzdneF+pC3ORw43KQaZ43pgHs9xC4TCO5E6VmB6n9LNw8sbH
a5GHmQ3BtwDy/lpxdG/q8CzUjtW+3PcwTm9XOVy5NPN+vAkpcD9Bcku0T1oHd0WmYAoxwYfYO8a9
nepFoSgK2TOcpYPWACUEvY8+1nBEYM/KL0bfPjCTHA7R6aRO6dqT4+UpTvrUwV4DtPN99pviK8S7
gbLODABkZPyi5+mT8kMVEgNhQBj8cfSt9JREeVEjmqlxXblDli1iBfCvaZVo2DuS5vPx4PcJrkc8
V7sG36fjCTi9499i9Z3Ok/O10KsK89j3vTt2x/EhUCf/ZI9fRuRBZkfEtwGN6AGwlfAbVw3K1JSt
2Hdy/zXL6tH5E369yuXrxhNPBRyShzSgnb2Br9Fv8GMdxWpOpteu1Spmsl+/r4JzDCw7rfVKfsu9
kmthkou5nsL/dmXmZNRsA0TbIC61bKev9iNbY1aSpbSAEVn1M71BKDCk7EQLcZjClv+Zx7U7FJKq
quVmP/CMrTLAqYREQCw4jL7/RBp0Jf7199jbZ+8ixecG1Nx6fCfd8Gj3SSle0fiLPbEVVmfbgABD
uukmiQTshKX493DnOY43CO8VtZMNobu8pqgE0xGedR2J1d5Y1dq7uzYV8yZdXaBHWWSHejvfXEIF
YMk1DLN6GkHrg6qq+ZkD9zoXrtT7rrksqn58cCk23CcfmOEJiGGMIV+KCJDWKuUwmjNxYG2bk9qe
vsipNaUn2fTjcR2V/T/1stzid1RJaMuMvRx7yU318rCfirfKJL/RTtp1crSHT0Hg/84rcyT2yTQA
nTkYHc5CSsoO2mBH8wnY/tIll7yoOm3AGKO3V+zjbyO4dJTKbKSLhitMIcyn4e4J+/Cop7lzOqbl
+T3DFEW2hPYJAc4It/tfy4hsRgSdzRHU5FqMQqZHEv91kJ5EkLxg7RjPmlZPqIWwFNPNMTVhXTlm
8KZf7Oz5b79C1NEdo+KMbVD0en0P7ZZ3x9j8yMHhZhE4ktpAp0hnyaxUt8b9d2rAD718+aq7Zr6G
QwmVl8lmJo84cYFNpqWfij4TvuwtW7GY60DF9q8IQFulo5BezTWxl6hcYN1OPY0qO4CQPdhZAVh9
yUXiRArxzi8zHEwunBGRRYXfRH+eLcP71xT4ihX+qJuSJ4zqlvGQaLZalAbKMLNfZwRAopeXrZix
xZS5iXLWGmFC3vxvemIoB5RqZ7qnJOvkLFF6lOVHHI5e5Qb3ZnPazQGUP9l4WCcjLJ9RIt0AvdbM
zlOH7urN6Ub9mIc5P5X0cma9Xb6kDtnXh5mUinD9PkhjsWbPImg5tE4tD+YHvuCCIPKcKMuF4K2W
zk8ckB+2kBOA9dVzXHnPDjm5CZCalbQX/LpBxewcqNdvNQG/vDIRNP5sfn5E64pKiGIWLE2glvCo
/lyYMG5tt29bh1KouLdrYrFPPHsrimnWgr77XDkl0bCB0ezREkMIYcawV9FKFc0i0L+aHD6CuiCj
BGv4KSiQFypxiCgn9fwl0jcsgI+dE3NGeM2I+pubfUkHGTyy+jXpCoa8KzPb7akA8XN0T3Fd3ilA
1qbDoNU30T6u8FnXOJ/j6T1al6xom8dK8XlSH3WgzUKMU4AelsHW5N5YSgIdRKf9aZlbr//IFOKb
EdG9QkcexTE6OWJe75TzWpZdam8wM6V8zvJbJ52XS+gtd/EEoGh3Dvg+JLP30RywW6a0QwdWtkIL
5ujcMc7yerRGgguZag83NHlt3F/L23VWIo7LyfGw0imw/VeOAxW+M+U083g5Kbvn0SnxDJl7Nica
F95tYeXjvnLZ7K98WlvsLEihRmpffGxor6o4tgpH9Zj7HzAZZZPLyVZ4De/DVQglVfMgLfURDDAU
xB+bwMaj1QoFqbmbDP2RwsVGpVSv2mm1ow5HrQ7+xJ/1mG1R9U+d2ISorhbnD9GpdHFjqdkWN5ah
3fvTRNfhPYeWf8o9EA3p1C0gbPz8/aREbuleBg3EqkyPq79wjp+qnU/8jzQK+byK+3cLPZWD24TZ
SwuS5msNoHGk0qyXFo+cRZD9rsliibb0WyjJvXbbolAmC4mD6wvwRdMQnorYKAjIh+HYDzg8+LwQ
N8Q5r3fr/TIVyRnkX+14WaV+e6lVYopwMWjNaSg4FRyzPiw0Nec9OFbQfMbNNaTjlo2sAc78AIwr
xQLtuMz6k/HMp4S16NrweTFBY3GzS2W9V1odFwZ0GN566DJe2CiV0+uJLw9vrnXQyomeac4MtAws
cRhetobTXDG/TyceFVvz+7zazjVPm104eXqpHVbVPpz41NBT/9Q2FQ7fJvFfwvOhe40UL8MBHG1k
POBNFyjgrwJa086OoZKbelbqHoGmNuDYFHV+cIqsN1DLOI8yiepUy31Ca6V8/zUjvQPSNONO5+jL
mBQEFDb+i8LY7qbKgytiNw2m31jUwHs3hhFrf7/DFW3VYz8C06MLc67yQY6rdjZmtv2R1H8/9R4t
v9bPYRd7zhbUpNjhcWnsGi3skedPz2NrongebuItRszRRC25AmgCzRdQrAkulXcE/6tlv3PrvYJL
7MDcC+ZYxnCxHsPWYWhWNzszz2ZpcDtrQjdFLfGDbNMVtv4zdpuWo8lDYDipBYJ08itxlrxiNRxf
mlKc4n4KwlFcoZnntgWnn3vC5ySQRupVncTVoTuhm8i8NsL6oy5ziwDCmHbhPm7/Z1fZDU8inKqu
3qipP57sixD7wXgMHSmUGM2bWNziDTICFKEo/8AJ1XxAlDmO3ndatQ/IoU885/ntL+mk96ciwms7
fkTDdrz7mNBohPt1IejD9DurfkuB6Wr6ZP6LU0rvun5FtE2aOcKZgx5nqYhL0U6a28tzlWe95vhd
WmkvcGB7wuXhiCAq9axE0E5O0kNB/lRje5C2QzoroVZAja9pnguTg7Y5SjQXcdAhIkPhM/di5tqO
ik34qo8JjssFq4yIqA0n2WObFaoVcAYrzLkRJI3VS56AWPeVVMOL2jgptPGQ4pat9FgDiI0Ujzzv
W0ygGK7Wi0inZWQgBra5CXDhOwQ0Q+6lJwTngGpuFeCKYZdZkuFlOciAGe7SNdilYMk/TvhjxFeq
oc99xRcZCe8/JNgHvzT75H7G1N4qoT03kjd95QH+Ijt+Qut8uQqQ0Ugq7PGa7xssyF7Kc6LffA1l
jVva2zNUcOss5YGd3ywLMDL7bGMQSYWdHDPDOHS0DPUnLgVxjq9kONt+XP0zx0jrr2aWIuCShRUi
J5/qKhXd+Zn5NQq6ZAEBYC6azWSUDPDau1jkmdOLVxa21UWBOdbopCpygMVtSdvbwgwX6uw+uNWS
7XFBB6GOXyrFUq66/2afsTqCY+/14dB0vVHy/7rmyuBPbxxyIeBSPOE4OOkVy/Da1u0BW6RPaeLx
EI/7PQia9vLlCist8Ryvaj5XoVY5T8kPD+HUF2Fc2yrcrFuFBLCXIf2XvP7D1XBoXkbuBoQuIGew
QOOU4XmRUW7itpMk+fGVp+DCmVOkw8DRDDCXlPg6Y1qd4n3Fds81w+9HebhjILB/+1VRgId+5VBk
vHZjstPc+KOGOYds/1MDp9DUkwfK4oCtECLCjbEg6o9AVaXyY8WoScNg/mr4T7Pw3GZmM51ymZv0
BrJ2wwiIdRUWocTlG5kQDoHux7NyrFVwpEE1nvCBjvhXT3PPZfEeW00J71wWUTBvGxWgxnf4Rz+R
5uLt7ejW6pwIDsjX8VHD/3ifmz+5yWRKfazLBFsam90ubpgYo8pAw/dmlSiThJ/0lun0xV+BbVji
9ajmoJjNJKcuA4tPUHg7Ejd73KINbGk5Sa0EEwBjbkPFYljdUt6o6yYdVedan/9BqzXydY53fx6P
wE0HO9Cqmgajezbp1zKB3hKZOHa0AeKf6imQSjtykP7zwJG/lsqDiZ+TbK2OOMjKag8lD0GG/hEz
k67JocV4gkQPKRz0AspTpg2ftRRt7r6LgfFZ1E0Curfp82EiV8E7Br8DSYkB4q/3yvBC2RAqEih/
55iAay37ugpRv0XwwFihD9gbb/zC8DSSSzejXR7vACJVrQlYvzQWAJLRAFieTnIHRDnwxkH+mFnp
+BpWY3lZxAvRguy8rK5vB9OF8VvdOHsd/x1ErsrwxCcndHbgXEDfqlMziuIhvH7bdOWhU1rSKXNZ
emGnQ4coMwCAGnj44JIAkiHeLle+k5nubIEbPidjTgam5FgeG+PmlzmkSKlw2+g/PIEupw+pPmIU
X4nnJlJkmxGqrEYSaaAm4XWbmn1Ao/mXgr63pvYydFwsrv3fS0gy3f505CqnzDcRWNP+/mp2E2Lc
1b5OYYdIpLF7iLWE08bbPSNGvRF1/8ZnOQ/tetOZHmoYfAwFHQMevmNt555mbSL2n1KLaDBm0OOq
DDUXt2RgE9Y6O8llbKuEWH5gGwekD0GB8NwQqqG5cor9B4dpCxGRgzkuezpWtpVdqYdxBNg90JG4
v8tIHimAIcPnH81RcmvAjDgrLz8uZge09/mHf/08beHQIRePElxGwyEPQtKhtsLYwla/T1XvCQ17
kBx905+5I6vhKltHlN0oe1uLp+zick/U9jn/au+rWFv5t9PsUjSzXbXxnHTj/kZD3Jo4S45NRfEw
TBSkL0t1gq/jbrkKwTUG0lEztHr7+or7P4Nhyk5qEBmaFB2m6/Uz27rytaxCT7Xp+JJ5DJjK/vcf
r3BLSVdqTZZa0LRUhlNzncKob5m/2+cZIhhPW7tWD5lL23DNpjHPgBrXbH5gq1nr1mJWXFBIOYcM
/WFPHC7Xw66WKtoj/YieAMn104IusajFJfRtjaIy1kAimm+EIlT0QKL/NkReuOofcFCAt0GFlfl3
gbQl9KQm/eqWXaMymMzgJ5vYI4iZwB49LgBzVhe3bqyfPl22Z7SrX3D/LfOs87U43pvjKcj5hOFs
keb7NbA5Fr5rn1+n5hIeBN89HwTp4GIxs+jmIGb3YPFPfigBfqT+3zIBUmVNvfQ6X4LnF4V9Kr8N
Oi0VsekRTT+1YyyvBuOLP62LyD8a57yXwmqP4K75QHjKL1j9DT0xGNPkOOmt553mBL0lRkDlp0iI
PjA5tlG1KBf0ZuH7GYBS/42uyK0L1S38X4ImEVp3oeA8dJNn9bZ7oJ/iHQugRPd6HCnVKP/cjt9t
hfygta08rnM1iVqBamlhxT+t7QvRV/+49J7rrG71iUmIUyUvKib6bHfnNQXEAHxOyd/CGfXcc+Da
LUxcEdfZ/T8m+Zlr3SB4SPTg4nd4tGkXGrGsonxry8jijikdEW4fr436X1UKs+a3htg7tHL2YmE1
RDctqPRQKbC5zF6Bg/dHHQvpVykMywBWdeLuLAAPgwFTrtl4dwewrPBRqI3fWVg4Zxj3qLCUuaSn
y1IDATwSyaqlAuTfWeFeItk+mR5VJg2UtvxV6az6lMSAyRIzlgnnf91/K60osbT8eKcjdyUXeNtd
8unjiTuafTuNhGDnmnY/GxEv/gWCUs+sjnS5a6NNuYXXEAdjuGO1TZ8ogIZkEVXyHs3yIGSLv0WW
ugfMt7vls3y4bSkUfkx3D1yzreW1GpUGeUoT7ACrRSYxRYr4lhKK5JzQYn7nJj9LOcMFL1bNKcqP
o8yk2Onie2FmEDsTl6Z+i5MDclH4SPmADwBbTLN1vcKsrvEt4rFdb5OIbG852KDlhcBfw5CAFQaT
waZm9ifuil3T53Cv+vEAy3tlue7IKa32cEHPzKU5fUydHaNrc7z/7wzc2pEA0ouD5m1tLwIm5u93
K1B9FZOjvuv+0uizvTW4pnlBOLvPoxfBnkVQymYxapLT9z1p1aErhGqFbMW/FzfoBaFAbYAZe8gr
zxL4z5vBoZdc/fttPM5YvXj//pICM3+5xAcP3MfKTKMw2fyzoJQi8QWecl6cgoUcSwJsO4RbuvFI
zEsHcdP0ActA6YIWUzprDs7bFeYIny5gYcijZWlBHCSZvOQmSWzk1GE0X6i6RhCQS1Zt3Kv8LhlU
nQzSe4AJ9Xn1ccwEEI5XQ36lLrQvfVrm9xoH+27i17e4F0brBCywJijRJZ1HcG2R2qNUJ2AUUG+T
6vpdTzFo52H1SbY88mbDjXNcAQ3Co2GNTP4j9M5w9kf/Fzt2qdUbo6APtlrHOpDxku7NXZk8i2lh
YSgHzUaykcvgJoqwhY7bkQXh5NUCzqTo5Qs8XdihBNGpd33iDtqqFpxIfolZ+ZuIdrL0sbcsPJf1
h/AsbwSMhSTajh8hAPb7NxEWFRG0ZoDqpdDsMOLdySva4QJlfwCN2bBsw63Eb5pV2v2huonGFqvg
9h9ccV3W3Qn8uS+ORq2MMPa0nhDNXlvqvSeEVWvzxPu07eeQd+qGOBJt0Cfc+DPyJPlAf2GXFyGT
ErabJWONyk6q/Oj7SZrS+fJDBd1sJXL3UUDmqaG2KSToUgKr8dOQBc+v9D6f+8UUXB/vd8ZjNC9Y
FySQWYd+BXUvSTeWtBxtlqXycxmV4vmg63i63rd66EXzd30PVUNvGbYLGkqIPzM+uvoLP2D+o0nW
3fU+TBfauMeWlDrtSXYcvSvKKTtwMPVubCgEdgOiOHaRJytDwEANCPIHwie1pLxr8gHfG2N7IQiW
GskieRFsm1dB8GXb5F7WgHqLDcRaLKBFysr9Htqs4gXdbHu5fOdUA7iTT0vcldp1D0xuULLGj7Nn
WjLN54qOwX1pjef5fGYpWaG5uvei7rMjFI6FthqS+bD/zTB/uC82Pk8yAbBGcXnLTviuf1PcfI90
Pf9YG2sYWrsZzvD4H41fN36Go62R6Yub4G6sVbuh+g/C+1DGXR+zI2389iDSEvNsvto3WbZWPj71
LbptArZyEr4g1m1sg3LikQl69TPEalm2N53An/hK7MOmz88g8m1DkbU3YOiWEa6s8EN+X5Z0wvTK
tSsSb+EywW3XyXW0onFcupZpJWmFRgyT04F192Pe/2mnh732HITeFd48O5m2uNf73+hSkZI2/jVl
rLNCf/XhUAH97+hCF2SMjr27ABwsDrlkJtbLgWOX8clPkFMiojWLjcbwc6HMRC84faFvuElRb2w9
xQJR8hHDo641st0kUllaZKwtesFh9/46l//lONj5XMZROu04iqt5e+9qOmp3MDzJKpNDooX9btrr
Wig/P3Flii4fctxgOKwZsan3Vx02h3vtJ/zLrFLJoMl9yw5Z/DGlkGa/VSv1v1M0rtQ3zWNCZ0mb
O43bsIOdPGUgQcOmwkpXIdUpEo4L+c0WoSGG07QzIiGaHKDAi6luD4BgR3VOmSH6J5vzoXONEizn
O8Q1gzmBE76zn9uN/tpqWeh8pNjCU50rKNJEFrXLw4p1xh/95JunHXDcIcvn3WRCQyUawnjpkla+
6iC57733wX9HKAOJZfoFKLd2L2K/K90ZCmym2XAwph4NMYXFikbXomxuz71oYiVd4t4vtq3IrSBv
TX6N5BmxcjcGwYYhWHrmvQGUFCLn95gwuRp0dJU8EZtQpFjWAF7yGTYNnmbmlTM7WT42d8athgOr
rW2zOLXF/vMlXMn8O3w+DmL4nYUh4vuXVP7bWTMj7QLAAmOgUpu8C2gnkB+/I4B9W3KLHjdqgZWv
Tu+U9UiKZtk3nHNVBOCGSd/zFX9IFys/KGil7Dyr4ypq3ayuUIJUTSoKZuOO+gdx986sUBfuD4/D
g2YuuiGLNagTgRkLCxAB1OceE4FukEqr18DHTcEKy2+3XaVMNLYsN3DNnsTiz0c+g2yTDZBxhYTd
T2wKUX86PBw1y57XeONnuw1GMFdy/hzV4TNI6gAmkDAQTo5vConVPfruMflh7m9ZD+o9gE1wrTeT
8AAK9Dse9Jwa8N0B3AlrUVx620b1Wqnuwsmna96fzbFun2aYbzin4zpzU3yD4yNG6Xxj5HfVg73b
8tf0KoP5J6mZV2DTIUQ52U3OZ7QvgQ0yOgO2H+SgDn4zTJ0FIzGaL9NArGMRyio3GZ2oaEFQXtwH
G0jrdoLJWH0/duDWkGkMRoWJRKdzuZBVilIfBq1uHB2c6q152E5Uw9DaOdKGOgnqoPVwa+FNFtma
4af+H+OQZXJUxbwW4EW9i+i98pGm1LbvCfUG5FECGM4Los+10c6QhP6tTmfcbVyTMWsfJHsB95mS
0mQD5ot/ZME8AVOBIyDm3dfrW/JM9vIUwYJQhW37d/jJIMbeIvKOx69YGhECXgiIHUz+N69Mb0mR
obWtYik9UfPCx19qwmzcvf5ULV+AuPpjre0kZyEbRExEITmMGadiOP3ZbJbDG2EhWGB0EJHqVT/1
bEsdFpemBRgqTrSfruU7ItRZQqeAG4Hnz+7l7szXZo/OARMXA2BmVIlr7lU75ikj/nFyqQgAKZQh
cH5OhBBS6Xr48TWqA5K6lHBEqOD5jQX+cijHPOkEM9pLtmlna+O72cF13Gn5hbNGSKaz25xhHO8l
qabD/U3+l2sisL5DuoA60bVWFDKaTCjfPhBw8WPIBfcWLKUVMXa7NDYdUjn5j8HRQAsCBQ4i5Q1B
WKHJFb6Kcfd4I2sqyojS9GN9UlWjWtPQW6d6Nv2JN3WELWbcX5zHOQa6i+Uuw18lVNjXZHAQxjMH
t8UI4fw9tR83LsfZSSCf68tIEl6ed0ujSnzEenZD97OVXqvIGM6pxuJo9TB6+PP1L8/x/a2DWl7V
ztSy/CA7JGG2JaPLX+vV5OpTMZ9kxOaQ1mxoerUBjWFGQnqzeXsNHTZndjGKoMWXO2YzeYZZfbXt
q4BFl4GknYaPzvpSzCet8QD1Di6O8TO6ohel9JpJ/mlwi0efIGgC8tyMR7hhE2r7G8F7dPfdt1wJ
3eI94hY2iheiWlxI7mmet7YUgMsZalJiJ5t9b2gnAZiCecaYeR25Rx4lam+k5zoy0r3X2M247GjB
G797fJlb350jqSwU3bUg4o+z1r7JlHGedaUBcyDtdSmPmyxEq2cFAqYIbYJxF6nVYIQd2aRT84I5
eQbD4n4+wKJN+QEoPZULCLk6mX7bHRhtcze5eY/R+LS+SIFmrO5vR0eUd85Y6kUJPSaMh8tFjv4c
Nd/CqzeC+WdodzTwFzZ9ErVNDOCQHJYIgEQeopKikNPWSo35+3K/UGIpOgDBZqyRnHNhkiFfAyxR
fCMHes2PoP4uKL0s8RrshD5Ga72NTqhQNWoan+Wjhs2+/k/oyJcUOvqUtHKrkUBKqJ5SOsWIE8Ei
5oNyZ7fKt1jhAEGmxFkB+xpJPo/tDMAPljif5TFu7rV0GfK3owUA0xkFF/x/VbBWBtBx0GQXpzJ7
uloxXT2O3vP+83hhBpX77F3PZOB104Kei7a40ytRZc+T97HDIEsxiM7+w+6nuWZyVFRDdUC1WzTQ
al89TPcxIrTwvDMn1CMX2+EfMVlMinHadX3fMV3swHJ1IPETARUmjs+IIZtICDadMY54mQ8wECjf
w/lIHl+z+YN5ajazhagPHe6DQ0KyDV7SOibfDkhlWOWG6CYo+DEGAl1bSR8qqKGi1r/yk3OvL8wW
SozPwXsxIXrmbqhs1YKkY+1PHW6jUhtTpYSR9V2lP0yA6hjF89V8USnu7j6azeoAHkg4guBnjOn7
U27nhYGomGh9Y3hGJC3HEz0dJkrZemPzvgQUw3ARC5khv3c3ylKNwD4SAuEG/BBqGyFvk6r62XEH
3kkqhj2ntmwVMqkzd3o2AiWEzqpNsCxdbU5Y666czivFYK38k/Rt5a/igSb1Ps0kG9zjzKwRs/Xs
CwzJ1xQm6srRqx6xeBHNrRiJBwz0I88R7xQ5dfrOzl2M0Lp1U6QAOKnfCZ1IsZ/vprnL9+aI9cpd
v3FN1YQriq7XqV/wkQLEeRwtoK46rtPHDCzXUqD05lHveJ6YY1dZwDg/YEe7pJF9bhzz+gZtGgKB
V03nNciH+W4wO9i7qYxAlU5w9Z34fqVn6DxURFDeqt8zzRmhW+zsFE26y3CU+pQdw1hY76AOOFri
Y8MEQHzfUVVGS3v/z0TKmZ3tX0QU4gE9leM8Vyt5V1GafS4XGOtOgRr1bZ12ofU+u55f+6ZQJmfR
4F6XqLC6imNj/xp19bLa9y8WMhQB1vxq9w8FjUDiSTSKjYv/I4s4Sj5CdWjUR8v+M4f/LOf1Z9ia
RVHo4lqgaXqRhyhDqhzVw5bA5JqwQwLJM+ENkqrnYCuyPHTEbfmurUEVHH3OPCRzxGFTPRWjsMBW
x33kgcYKcxEfTPTr5KUCETvLgLh6jI/BvHjXDnPDZCVB208cWEGhx/QplKYzbiG8+BEQ1H9Tsvj4
dNQ6r2gqxzSw5xCTxutQX6p3/KpeNDHNez6L7TE4PBBgY0mGPQjo1PIyeWRK+nqUuU+IHk2r4O1z
Lh67g4gkiHoaL6Sz0tZx4TXenVOZ8DmOwz/5gdAmZHNIJvBg0tH87Y72b49XVuFHKrvOsNT6M8xp
mrLx3bdwZnOCbKtTrsbGsOKAmfKffP0fRwTApY9hAfhqkpx5ruSWGJ4WJEabVOS97vmMkRRRsJhI
fH5bd2SHpQMHH2fljuJH7vW7L+8S2JbijOInxetnzsgm6zfoFkL0zji/ANCEFp0V9RRsf4ad6mcd
N3ASIPDMllHwBYi82MuI9i9cPXuMnniig5LpRE/d/Utq/OTDQ+5piePKrmkNeygKOhsexms1zWd4
2sUeJK/gipzWmPKa72F/6/t6cXMOT4CX8PgO4Rh99AifA1tOOo4ZtyuYRIZLZkMXd6VRMt73wl1Q
Movn8RsoyQh+9GCf5Ql6l/GSMA3KnPS324jmwruy28puE2CK3svHxm6GujCCkfuMi9PpC2x3T45u
/FbZUXaSRck2Ur+1npP8wOagwSx4HI1HuBbHJqCAWaXBVFxjLLmge4RHcuRYjWPr1bK10KkA/9pf
uYffmq7SC37fEN/+Mpq7I1T1NeYK1B6TO+5682tZuRSjH2QGP5zPbTmSjbk2/MqMjNSTEMAqIeW+
+Q/uxPEhnzDN0sFWauS0FtluKBvsrjqBsYfAkDVn8jlXVgt0QtxzKWAM5ll8O46WPIQEtejWuAIh
s8j16usUnTgKX1PdWZG/jIqKmw+rVc3SN6Azajvz4OXnV8EjQAS6DZaCN29YVANxDulZUQ8rCbNS
kdDrbWXIfwseWg08yhvKAPWsjO+C8RF4dh6XfcuzZPmzewQ71Yr2KAuOKkGv4rhWhgK9eRwW5gg2
Ky4S2tc3e/UiRo4lMkoqYaEK2XWNfTRNqGjsthOPpk3hhc14OYibWYyXJQ9fWQH8Ya6Vugv4ofU6
gmYl1iWPwLA81Zug/ftnSrlMb2NSaLdG6eSr1f1qeYitClxrT7c64lW7C5MTKr5ebO9dcM81Y5JU
fxRdxKKqRdkiA5wNkwAmZLznY7KjMWAWMp4MxacQXtg84jpwwSGkz7kanW0hRvEejAPt21t6OYc6
q/Twh7ZU6yrQOlF9EP5fTE5pgi1M9mkklTxVQig9OxIPcaGyKRIev1sv8yjKAdAqLjKhKlmteSUO
8xxeih5O+0o3xMgy2UWw61cVeZPl/2XIuJ87F+m51ZvmElsc4nb4ROUeghHq1ngF7xP+x2zddTOx
vCJd5glcoKJWCcTyoDz6pVdAiRqIRAZ3e/MF1STea2VxZM9O0zT2B1gp9mdvxveAI3JloQlAWImm
++6bwKwHdP7nonGZa2anL0AdNXnobZfbnDwRKJltSu3ycXUnTE8Il385SLJGFyGtUTpAkOdWSBUB
lmA7d1z8uao5TQuMymXpGA/I/vho1qKwrhcXx2SK1DQTT4t1FMYs8GboFsnCXsTC8hOwbwso96O4
McPavrzWpLETWb4UlBswz2m1zksB59rz7lJ5uuR/XUV7BPRa7wd4vyM2N2iO1lwda0OLbtuuRR6n
yK/TEpQmpm41TaQJQZGpUFpE63NokMPHLb6UTyNCCgTis4/NJTAbh31wm/meUoIAFlx/02Iflwyj
YCZIbYtfxBl1gsgmDwxdxC/4qFlI2Erq0OlR9vmj3XlmEL25uqqXI+w635mv3+LtLZn5R0c8jVQB
klLF8TYK6ivJk7MLboMCYlpoWa1c5snobMBIPwp5tWiUFVTp1bewhGYxiICQFjm12mDFw6DScimd
qjFjLWEu+HNkdt+W9i70mFFpIy1lKA2WdUWeE5XUgE2Y/D2+Q8FgUSjYDbBvWLJ6hn9WYsv3lm3V
I3LIowdGVnWBl355+9liSHQK7TvQ0ODpmTRHXXxtI+w/DPvjK7KzZ4cBpKVSIJ/dAxRtXYgwWuTO
2Ny2G4btZp4ywZk+/0uryZVlqE3G+jzAKYgvTAK0o/iXIt2QGbdKxJADHrT1MCPxRroB/nJ3CKvd
w2nIEqbfqObQ4NP1wJ4zGSANlI6AWCr3MJMyVZioIwCPdRpf+7fsYWz0iox93lhVOYk51YS9MucJ
Sl0kR247jGhQMjGpYaiHujKNQ6xvCVa/x7hrFV3T5NOxMtNkxiqzBYDXXdapnrq/SNa6oYN4HtbZ
II9tWgTXCnHYAXGRsv/On5QbJrN7vxAZlaTWPc8lbgJh8uU8ZZpS/k2bM588Gr+svf1MmCPNLe+9
6eBS+S+ujTmHTcO9WLE2RF7lU/JsmfQ9jJKT6r22R4gaRD1xqphJEU0mPYePTXaT8OSU5+pFxxs+
vNslB+Vzdqsa3Wpq2qFkMpakV/qLOHDD2DcP4wPk5CWXllXaTJL0mjPDZ3ztTeLwvZ/abJ5wU5dO
fhQn3edIxrkiDQNHGnlEuawXEViB5oAnZsyq6Bu8xQhN+pM24Bjbmf60oot8u1lWX5uVqn+c+d8m
nb98I5p+Pad5jfQX/KJa36L+GtKFDHmibWMuH+dwb7NVl/8enAQxKEYjQHVjCslBFAxcFUlFnXrQ
NlH0CvMQJrG0I2hjDSKSI+dHyszag62hk8otojhthLZj89crIvyo3txindNnVBH2aqTj+nnfTMfv
3OXg6SF91gwJBEmsvNIsCZiBnUbPK57naKyuutOtz3FH5w8jCr11WM2GidFnVOkEIjU3mdZJwFnB
kpBQjx4GA+MMKSKLe1XNFo/fvn+3KktzStVpCeiXwTyT7x6I/jJ7Ie+1hkHDIriu0K3ZqzKWKM0T
QXI6f4M1XESeta5dUw4HAPvA+1NprQoAx5UF4lG3/Ok/YUQQI4swKnekhBjqNiLtHF5mI/mx2k+R
0NslcNh/AjLwwdzgShkUhqDB38A+T4b6xLICZ5fEh19NcwR/RfEC08jnxzSkmvRnLTuR2jIrnTm1
ZkcUsYtDck1QL6rYYzuz8GKGP2dBus/a4JZXpLEg9oGTIt3BYw3lkxJ+hvyx0Q9O7EbeCGPCu9DC
GcLkyh3IY8fNlnJmMYCYA3vzI3Qq2LyWV0JZ7X/Znzl/Nn5SUit1MPq29b00eD2SMjYiKvOrYV6j
Rjj+YJ/ohlJaB3WWFfoSReLbuAp97m8CuQ4FrMDKtE0NqVBpi9eXkMDiNSSkpsFn7CWKl2NfX5TW
mPXtr+GNuX3Bb1VinB6LmsfUMiOR7jzH06wPDmKgk7YCdD6+1o1XMxNOufq1HWZ5Mi8ORdtH9FCJ
p7lDJysUqitegzG+Sf7MKsuplguXZWid/Rh+0dBBDVF9VA8dzLR6tUvpzIBGXW1eQYMV3lCotfXP
hN8fK7TPIekUziqHIWBdFR8hv8x3FZWOdQ0MaisbxCJKYzavkWrkQdSDWmFxdean0tNw9C/jY6y3
Ncm0Oi7J6eSYmuyuGaji8edwvpxEraI9zsw71opcOooE0OnaCUqV00Su5KQ5q0zKxXTRFgARVUdN
iW46VPpvBWWYGmAj0oY9jd+da3YWGqGmZogWrzSAfvG1TgycIy4tw7TEd0WrDq9oAqKLqX2m4yTs
M0MbcQxcv0TyoNZutDbRtzWIVohENCT2DFYhhSX83KcQQD/IGRDgpUW0pcOpj0A8Pz6flctbgske
NHdTpsIgTmT7b3HSfif+1wzIhzSG/FLkIYRbv9BYljozoWho/fzZpljJznmg5BxvW2Gy8W2twCQJ
EK82jKmbIzp3HA7uxGUEbvvM0G6+ADnPztguQl/vS1WTRuMSTAK8MkJJJQVbGoV+xb+c3KdJMJmc
ae59RxGeb76Kfpm7geix9e1FdkWvbriiK1O3+oTKPzxK4faEjpIuaSDPs/R5H3yYohXKHm1bVE5D
8wzcUdMW7otX3cUvykz9ckRz7it4HCJ/cpIlpEq3gDl8vr5MFGx/AXwUfw3QTXSk51VkhsJ3efo9
i/VMINa/av97Mw4dPYbgQLeQx8dJHcQlimTPM8reL2vqaDi9H5HYqAmxfzDGIAJ0p47LRu99108P
oy1LP7OeKvCsNf1raJwGmYla/+cLp3w0qbnTziBvQEkjUiDH4c7y5nHZpcHnxI4ZslF9YJVrvUVe
cp84tZuLwBeT/08K9IBC7H8trYBCQ6FUQ0hxMTBKhlumfNfLXszlPTEzS8yVn8kJ70qP96N47Eqm
k8iWZPfWj9XMQjOtpN4hMFTxDrZPLrZXgqqe276XYAoFY9bEwBpvkxYKOYeIoVF4HfYOSwWUXrn5
k5NE5n1+N7iMbN9Po30PBuHuxAy7ZM6uCY1lBE9pedTilfKW/gXyeXMw2p8bz0bpQ63VhQ38eZUf
HwBv0yKPx+UKD++FaU+aeuOGkoulpRJLAihTtmmpghK4VGVS95TKBUMyceq5KriRybGZIzi1T3rg
M8Z3S4oqe7qaVez40q/C3aKRC+beU9eLRtl03Vlz/TNOJbSz7QE7JcLxopVCo7a99Y5axz0VzeY0
CCwz4B1DZia/aSlwVECJd6J0l5LEL+gOPVsXQKhDIxXzC9CSaBcpKqgPgiAse7LaRoXEWJ5CWIJN
wbvaOQKz3ANOe8mwiLzAa3b0UbAuFjRPYAA8oFnP+qbZVZqI0w00WOLgr3vpjlukl0fFuZDdP89S
3QUARMke8v8VZCYGXoavP7bjCg8H+TFoEWmy/NdWsiQigWACf9nJ1szrIJN5LEKKi4nS8s1P7ni/
DHP1iERcZgmnubGt+wqdH2eCC23HsFOZzCGDN92AeazFXDm5CnhYbQFFKIQPBsr9/fQ9I3TOup2n
JaEZK3zdgR4l9RdZMA2OUbSwfffbp3zWNC4hnWXQ3LCzudghMtExkGGrI1hwnUpcQSgCjK3IDwYp
3TjSxKwrGB2/VYsRYZ62aO4sns7STlE5wLPzzkjiVrHW94SDwSPkmxc/zkb1Ti/uOqLNiO/ZQ4nE
tAOs5piJJXwsjzZhbC/WtkakhunwpBEm4dr8ynB6JmZXvgWlIiLr8GbNGq/mguevWgQrnGyzYjeI
/T3UIcgckcUL9JZ1L6QmPaM0R6bWcPlkhXXPhf8yAeCe7ROgxO96wLmCnhFO1NDhLQujMK4alreX
ACy8jgHxRtl3LzOjs115ir+Gsr0BBQwqkbQCytL3wYKQ2rFAcFqAxOzYbndzxet0tryitVHzMtTX
95QNIGesm1WywGcYpucWPyOGpkwIAEdOe65L8Zt6smUc33sQbE5vPaajRVYlFdA3AbpE5Y2VhfH3
BvzRfwHyyQ0vxsa/YR90vfAXFK8EO3TjD8GvJF9zzt3qQGwc1xxsA0v75uSth2FDaLPCvNrH8MAj
LnTfWbn6Bhe3ve5BTbCJSZBBV0LMj21hFUs2dTwgtCbEsX/QglQdlkHTDtu553f3CyxccqNPnw0a
VZO16qSR8k9G+acTa1C0LkmnaUguH43GJ5X47CRb+G6uiwK9rS8hDhEYUrxIsx82o4/TBUaPBAlU
tkMIGlxEXNnR1+IGDhRqvMVNv8W9X8lUrek+4nXZbu4SxB+sU0dh5rjOhrPALQLCvbwRcRKmhrLN
gvgfyuAh5vVLMA2FLE5xmjV95Kj5XSzTnrYnmshC2QsiBujmEiAPzkAvcdrhjaXyGmIPfiZ2M/En
1YCQF9NeJkZwCOpx9/nIFwCohhbZEzAOxMFPnNFemOiJ6SKMBlcWvXMXbWYr5cd09j1rcEaYT4KH
TsN0UDjjGGpQydEiWHcPs0AfnLFjOXQNtXsAiheLjlQkbjH78UFNLpDKRI7oCyZZEegzJKKo7igF
IGwCj8QsdfU3hR6cPhuXA9DenNJTMwmnH9MWYtwCxUCA6pQsjkQzm76aPttJfmibcvNosR9ZDLaR
TOu94uwu0abeSMh1FjrM4bYD3NIdgZ2J/W8Nhde4vPMuS1/APOe2CX4Pl5ENGZQ5EEin178FYOGz
x8wMbfKZHU+Yx6w/aF2qMtqNW7Y4yj9faY4ghpDugAMotRmGHTfHbULRFCABrr7cNe5DSQIEE8uY
ni1OJKBF+wSk1npcIhcmcn9SGu4GpSweNHahezN9A3A0rOGxzHT69Qf6QaJo95v+4MlVuwfPc3OP
Hgi+d4KTSTmLUsilOBLi51GWh/6AKHe9nDXhwvltbYAki9XTnxPjMJ5H7dHGAgG+1m8K3NVJdNDF
oh1HW2WQlF03IwGhE7JtkJifvXWGBxf0cXEuw8u75zUg3Bh19rSkzKkaMQnT8+D/zqrsAA60Dk4i
cyARTYbXj54idImA4/c3iP8kzhlGGfgZJTSkbYlBTQSbA016BSWTdFFQWFCyxCDA+hzK8dJODBjF
fxejxH0qrjsN+DvdTpNUQZNCuqudmehdokISm6JNk/hJr6mA+CLBEo75Qf7JETOsE3GxocTo2shl
8BAfwnqDjvfauyRMn4qB/2fGMV5EvDKRsHaWvnylET4p5X/daghxEKjlo35tr3+/ddDomu9JGZEv
nrdIUrHEqy2bsRY/TUEGAvS2ZD1arXIIWRjc14bvPdIK96+ZuRpdiTDX8KwFSrn3xAxa52A6+U64
D8Ol0fghR1hGkCTKD+R2yI9JTrh+IsR5TxM2itiBuGVDOwTvKra5+Df53MWwNuXPt+0xFTBsUYYG
m1r6V4N35ES2Ixg4Fgn6EY+tGPls33kAh7IDx6yl/aGCwzr1Wmc46cThBibjUIt8II1svC6uzKDQ
38sYZxh61TZYZQyB/yoRlADeKUfGiaEuyYvbbuZOZls8UFY6bflIpVB9lP2l4a9LVn7D9Coz7oHt
Zq7SnRFkZam1UAVY24UlDxkBLK9DKcHq9T/YVnGDqHsl/mQ0fp41d3pB0kc+LtwnLEWXTt/1Pyjn
M7sXAqZN3nY/5LMH7tQkAnHlTDjH8QEiWs5JHCAnv08u0omZwnFRYgDeDZ1INqFQC/3Z0VWnBbqc
3Rqwr2Hyh9ecdXTkiViruBwa+4OQ4a2TT+9Sl6TnqoFAP00ayldiSPOsAzm93k6hxzvXTsgVWlgC
sCOlVddPIewPpU0zw9DvZKeJNB/MXSBqBP4FKt3FkMPVymeePVhcABzZSTgswaWufjuJGanvrbxl
tub35dZTwDOLc9kgPZsaVZTuMb0zWXs7rXsORL30+ezcR8cqLw2Yx6QAMVj/P9TjLBdvGzl69I6X
9oCtlIR8i+0+klKYxz2+9rI5QZIu+Y0hKeA16cFHz2u7RE8IN54vPV6Ug9geErQ6oVlzUQsAtIFu
qCeaqND1GqWKhyHSV0NU4J9ztvPTS3E19/PfVysgx/NDFz3o0x0CVVcP1mlseYnoHpln2jSN0Rh8
f/1xodYOfH37ClBD3SEzGFSjTSZlh8NCMQIqG2dUhfS2jvHNIsKw/gXwt7ai2ggvgONnhsMVJq5T
j8A4sJd3W+zz+Ak2yptXMR288zN0MX8zjENx3SObSrcZoZAxIyQZv5NRGGtbd4gDolqg3zuh1j4K
IX+TbOEj28+s2iTKWMh/np/BJoLmkQm5XA4pwgxD9+Fqnz2YnCp+suRtSzGz/T8O/ONlpcEehVer
RXbv/WYAuZlv7GoMkxQrh32XTth//rdr0vRubEmRNJYz4VuyY0yeWF4jsydyQ78gJvhWLiphymat
GvmcLfbr9taOJdOfzwMZngLHExFLujl8ANpTjhKn81Qn/ED+uEfkEcWe2YcjGgCOutyDtzkuZqO1
A15c1vTPwd7JQvoYVcliOGyYHVvVe3q1VriEuKSBWcbywWAg+YSoWyqmkSwQKJ5wdjvS4LkpLeGl
ZKO6IDkYFnOsRyCTT4z1EZ7kKR4nLUC7yn4+xrbsVlpUf3PIOdtkEMR3CXW0g0VITWHv9LOx/7M6
S8I6c6tzD5OyqMC8NLWBLk0pSb6MCXxQa7uXgQcmGezKhk1RXSyOKjIoc7sUXHLba9s4OTB5Kw4R
PPp3J/6m0lvGug806T02motIsZWy19bQkbW0GprjvO7oBWREuNPJadW6VRSAjCWqgi5dRGwuOrHN
EVxAJ98bj4nnmKYeRXclcwhYYwtMiZsfm7F8Hx1j5+U3VpP81iLbUcTl+9q1m5K7n0R2lFD4SSYV
Z+vZqUkQxMtx6fuAGI9/+RrRKaAX7JaFCf9MNFQr7/TuvCEbE72qO01mGLjCbTLjV25j7QUiZTxS
zCfnQ0Wv4+k2vSrnlTg1n3tOUDo3Y7yXjtfAhzBEIggrjxJdVu+hJy4WWo4Nc1npRHocn8tC22Q3
JoWpkQUR9khxxAIUrd8JB3N2jggu/Vo4YGRvmRcnpvIJzKQyaIOg5aw2F2hjTkR+OwijhqFAkf/r
z8E0usFgObT22NXG84kdY7N65XnpU5VQi51zxI4cMrsJ4OY9aHt5wg0qUGbn5AhBBQCG2wp51Gtn
Pr8+zfr5QCqepvsy/ntn0qv2fqNtmwUpX2gFtcvt6IRUrtNE6a+VzzcJR13e6hsdUHi2NwNF5JwW
d4f/DSqGcd/tmoMQuV6WJ2uEP9qhY1/qHPUwLILUlN8iLZJUCyGt1n/MOre2UlLOaXHFmFY9KNDu
r+waYSDq8Qu5VgJCRI9BTPNhPN+F58zTWvsFNZ+hrU1kkedq/De+lWHiuYw7i8xybXZCvvzogGUk
EfDrW6JCNhHlDTzimV7Uy8Ag5x8xeecIN/W18F2TBW4AP7m25URk2q4BzpfaU681eO49Op+IBu0y
AKFXnmFprvrH6h3B2bZrWva4BxNtwZ+Tc0gznUdiu2J9gX9/4y+p/2hA9KRMZ23e7xLJcYywzrpG
4loJ0PM3Rrjcg2bKtG49AY8n/6UlPpn39YmIu6N8QEtTqJWRBmd7q0Pvo0mPoijfLo6L3aD6cvpd
yL8x08c3tXOf9jr5x4ybn9xgvO3uyTXzZHHVtewqN6NzYvPiWWL1UNmcu+mbc3XxBkRDnestYhmQ
2Dewwe6e7rC5yAxUh6eNhi9LEyoND9tsQHsDeZQEDueS5Ms9XrdoHwI2WV6k0STzROFFqBfLVpet
Zb0r7+WWAvsZh+/pzgAKiPn3g0A+J9AWVPf16Bd0UMV9gHGJhzQL4gZDpIX44/pM2+oBzzhBJAvS
DcJXO7n90DMoEY2iOOVTYCdgsif8efCz3lWHRtH91LSA7h2w08oPg7I6wsgtcqf8LOC4bo1H1eGS
NfmVXa9N8S0ssmt1N8Dl2/m2H1uE2n7cQEGJlPQwInCvoTO/81bTnUdcyLI9cPNHmGF28OUeUZAd
ZP+gaKD+esrR77Bq14tJ+JC8+1hTVMnmciIHNvtqMvbNLyhTQughxpcAuPBFj2JcKsxXH8q/awjh
yM+hvrzsZ3jxeZwKXqHMifMt6ds+Xo0iMXeh0si1Yh8cz38d3k03Gd/P9kKZaZUmSAI5Rydvvthv
s9iMgm/urTcwu0xFwuZdZmcY5yFgCbodXCotnnlWpLsEBPLG2S/c9CXpeX9D5rIxWx2rdiAOL5Us
trMdUpMebWw9iJSmPa3Qa9biAg16G+YyFLL8EvB+KFUeTM4w7J5uTR260J1cvaN21QBeJN4MEcE/
bb0CS9r2S+dumxDzwlTpPfCaOBIk/Tn0LikaLQTp2hDaRAxIJBkRG82ezFWTbI7B92SCH5kvDCSn
qOgidiM1N8OyARLrPVpozbUhSyh1u8G7ZYrtNt2NvLklFJ5mUlJ35/LsaJf8WIGvTwTL2KE8WgFR
kD+2C+l/c/kY7NMwX33mbgkVU8t0wF4NS9KfByopPcCOCwqK21gE4SOsvNVck3yCsAjq8ubV8yp+
ExHXeC9fkKcob6PJW6yUt+Q9Gwz04S2kXcQLwnAxVMlOi9DXJ2S7Kyl9lIstEbMNotbkIc8mYfP2
/2P0AiIK68pjcBiK9WTTcrjndCD4canlTlTWTa2DO6BUv+/h028CnAzzNktNiHNlyx4sHpn8NYk5
+8NGXwag0AI9S6Hbe3gHxBrkl+6DrcCcdbOTrW2ZeBXwPRVsAW4nK0SJMJ+xBsEp4DROfriJysCq
dKRXwIdX9Y7FGEJzY5i3ebdXF9aghjTXKPhOMJxX0gY/fGwRxObaYg7BsPbNYa1fAME7MsM3wkX9
+RbehXWis+AIglW6UOvEq3MAJIBjaZfxaEGRqRexhht26C+g0xRt3Bc7MCkOSkoER910Y4vnsVuv
B1y6s2ByUqDU7Py4Lu1Ki6zpFpc/sBaNzqTnO1ExsnPuCwtyvvzyMlk5sT1v1FA08K/6OaAiO5Nz
wY97W05NER4FPnCVWHZBV8Bax9KL6bqk/hv8UxPe2GEyL6eOr03qMU69/fKYH1C4gJJJPlsmXrhY
Iq4MRirMpCEJlAb1xB7jabVFR4/nO8m+2F2U4vlRJIlsnVvUo06uaImI42ScIY4JrrJOELDZd2lN
0esYMg5WYQNMJieHDE+OAO8yifs2e0vJ+YzpOhUUZbFTO0PgCT4B7l63qLMHuzrTYzMH35oQh8EO
k/CD9HVyOgSgrtQ11FwHaCdjlWbVu62FNr+AlgltYN2AV0zD53UZkauo/DRvmDTZFam3W4EHCIHe
glWOhDXBN2+PWHuvc/fZzRvqV88bjCrcxY5JCJDVfGjibDwuL5pQsqujJPXvIaATeFQ43fV2FrCF
whCICodilXfJQvJTZlU5sqxEzUW7BPGvMPDGZqxZHRRYF1o7Prd/Wkbz+g/bfyxzzp2Ygb0NCALA
OqQWf2V/tUHOaesDjXQ8mQuWRSYBEYJG8L7ymyON6zBAsrpjUNAA2XIEzwrOXPCMTYo26juehNvA
BQwhg8eEWt4p/BgpoXqqEX5BoY+LnkDds7CVj6JjTCOun0tLQvr1fh7By20/3BG9vuoy7QBKbyN8
8JvnJt/yfiisGYX/wl27ytsL/GqDSYobtKr2dYEddfCuiLJgnagot7aeiX6gq6smW7yPEPhaXmO3
Z2c8nsI87j/7DvJBT02UMKQ+xNtogoSw4ct7hnWPMlvRY8FBBoqwbD+tC2AqAeH9i6x0iUJWgR/f
+VbZqQzjnD3suaJPoNJHYrggi1ywAtX/zb249IUOem8SWv85kLPQmFyQBjdgjHY/Uk7WMUEkNBFD
CjPqXSl8k4wm0f+F3J3c+HJ3NZ1bRFwkTwb193kfXNnEW/Nwlc1UIeJf0wqNWq5Xpdb7wZri7vPx
pc+Y4UQ5yOgXjWHxUt6j+/7atody6feCsotn0UXYYwqa8iZ/iCCSgCoXUZKK7a05vi3RCw9vWtLy
rviFZUvGAfuHTMsmSth3Hpf/7phm+ItxZENqmq3z1VFLQBf1vonxli+Msyr+9NbYPZcJ6SDUKhgs
OnZYBFpcmpaxznouWQq7AXdLSQ0YdOBLc0VvhvIa0s+zGduprpFzzpY9QdcqxsfaJVx44srkG2dy
P9SJLlEveFrWKUmQFI4070LEJ104guKXUURXrvWat2+dgHDC5RzxnM6XvaqZxv6LJern9jGTud0e
vv9ONTPKX3ZrGmmZR2UV4m/D0q29HN+Z22smPhcfWX90kjOZvzjQBXAgLzkwWsCIWWw5c9Hb2ygM
6J/xPzM5RwhgjABG0edjuYOe/O8ClwvLtGbYXna5ZCu73AoePpp0q37H4EsjovgY8gi2NJVKuHUv
Wlo9p1u73zRSBJQvkyZ8SdGA56BrWfAXPNQhwgsTsq2h5ZUnz4OoHPuSMaG4YrKsLw2VL6MlRpPJ
R7CJ6aGmKJ8HfKrFopfItyHcm59gKB248jkqrmdzXA5MBJ58zc2iDwYg3q5PnZQJoufP/qupIxej
AqInJw8inKHdWLCz7GNDqC6kv0lUpJP02jJgmW31cdiq8ebN3gp2W08tP3G+SXJPzj0gpfH64Tr6
/6mVwa7qoE2NdpkiDFO/oVqCjjuEKBMJ7Ku04XPmZlypyoK2k492yZ83ksWrzkTFRLV+ofN12v2o
PGjUdF2Lt3kg3GkPBCkQdYlU4MB76+YdIQaFHJAbc3+W8usdrCNx3z30NDLSsDt6r7IjO2afpuyK
ezSsCoCP2eoExgE9ViViCXJtjMmYWp3yPshfzWbS81nbu5m7zDLMBDNRXunj4pbvR2a1APGwUlEA
bWFtN9XfIn+VSqS8wijZ5ELAXUJk/WG5iQRER2WYVXiBgVDvRyLJLIHasCPoWglH9MfiphmsuLW2
ZTwdkAPLOIo0sk2sJUiLWcRxj/aRtaqrCOa/r0G9L1bn8o8TroeoN5SfIOZ5Fl6l12hMjJ+HBbZV
7E0a24EIJ/eSRZFbXkca8kBdcggmMyAdm9YfWLOCy46crbaVOR4a7NCOnyzVTtxtizcxIntvgrUY
zkQ4TIqgVcGjMXlWo47ryb3Mbs4AyoWz5hKSt1lOPm7cZFtvTJ8f5YZ9p+OL/vncMu1PJCsLnfSP
0KP1KgWaQqasUji82X2A6B33bEjzSUnAkJ6BxSvrwsy2kXY8eJ2De0youP+0f2Ejm8dIJTIgb8IX
OBWkWMr/2h3SRlEzLRaUa6SblpFuWRELscjiy1/e2yc4KdJQOtuvNcvy0NBHcgmQr/89f5CnEJrW
3Nj0fOhxYutBufmtNPBvmRzBK4opTCHe4bFJJydjRmEfLjeMuGYi7H1Xe+HPCVacYn7fW1M+2VnJ
9t2GFXt146/K3KrJHGFxXVOqVtDAqQXnyB+TgP2Aj5i7a8b9Ag1c0Q5zPCDee5M0awwfrBfqZIBM
qL9cc2ZbXTjvCWsbi+Q6BHCmIQRpuLe/Ibdaqr40q8ZJsA6LU9lcSt4aPbSP8LDLUip+Ln4O+AgG
OIA0Hs7lffB0azN66m3q4irkp74czyyj5qY1bS/4gX2CTwlwBDEHLFNQz8tgQiSzcw/5g1pGdrVt
Y+N3ZC8yN90vJ8WANzKfZtMvbX2JUNK8+QejvdZ2MZPYbZiVNkwtLOKo/0vsPXIa6IvofiuS2kBQ
DgpqNqorYaqbN3PXWipwHCUslKEvSuQJ/+hqx6SC5Ab1gAodwUkW13+fO42IXBFfdMgItkjYmu5s
zQw3bZ4a0V7dRJBiHWeB5x2Wm2FbNL3WsggFlHtrMBDom4bnqggwPBG1JVSDykiEN+W+ed0F+Wym
syCwMvaAhZirGWJmV+b8M2xp59r9qW+4s6zZzzUlPKWP2TR1DMibYu2Im+iX3oZQKVkkjyvmBeFR
0xlSkXzYvmG+CPQbkmxtt6g/tN5SJT+r7rYnGPFtVj9ZiPnQOQ0Kfftzt/xcLDPiWSecYdOmpHZw
IrF/GvEUo5seT4lGkQZBi2J6ZrYeI3w8nhgeWkiHMLLrxOSCk5+NuwBfPVFMP6FwJae8cI5TDfh3
8mts61BsuVi8vmPvSgfdLEUCGe30MJcHSApW66DxIb2ldShTsc5p2UWmP0e8EABd6zcwfpXLKULI
D6xT+RVyT22krddxGsZE0/vREGCVQij/zqPMRKKzqINMoSlIl2EbrcNiK55+sT3I0jrX8G0zwDlQ
jcN0LbQyNg4cciCLGweskudiQGTnAtnJJScyjwn2kn1iLZRRfbZ3gViqohUpABmhlXFBST/UKw6+
58u6oo+rOcNdjD/b4d+kgMTWC6xF/i5r1K1fA9nES/+YMph0qgiZcwOGoGf66zzBskhB0Ogxehos
ZR+29K2k4oOV+QUYFDS0RJ72732FKRUXR1+E6FEB+fwnUrrD0OdlTvMK5eW/APD3ijnTa9uPLU9G
52O0E8JC535u+XtFve23ptTlOZCOpPTE7PxpOog9at79a3Hsgpvl9iD7DUr6K83AD2mI4ACsiNNa
W+uaoH1ceFJdIQ+lKJcsf6AXYtfRGv56tchNTYv/rljHIBESEEgJqRw3V48H3vTZfXPxoNJQJzDJ
UhZLiKmjsA0YsGjJ62OZrWLbN9l3mi6vsY6YCqcHPuWdy6Rajhi6BV2+s1ErQ+/fK+jmHs849gBw
m0FUn8GKgecXGQo02Ko6L5Lf7f/a9wJ6us+bf8VBLUokXb9NddbdCH8Wz3qIMKUZeDDMXy6ik7Tr
/A3P6iaHLef2m0+0EcCy8HGFgxpfs+cp05bmiVxrpkyI8rDSvCepmBcMyBdnHQWe1UnykRwqJRmY
dIVbAcSLQtnzAo1+gl06f5C7RZAY9duoBDlEKH+/rT7Um26FWT3sa/RTvOFh8JYpeoW9O5qrOF+z
OPJ+xZOYS+YKvorNs4F2AFGJRGjqbNfGAdbwGXNGinUazoB40XA8N1UjQVcJJ8fRIHlukFp20uoQ
whduVEkhoAxAhybiuGnEtfBGPqgGMkvaViaTocZ77sjwC1K1HluOjOQoD2Le/L9zmE8a4YHqXp+T
xfxYkXInFZrcSOjrmZUj7M44mnEudKRDhHCSvWGStTVkT2QIx/vU9eQJKmJFfQ83KkBbv9zjYvR/
7RMoXYHUqBzstVBZvVfluVkqQChgIdx/AJemvmPpFA1IiQw5Wkuadd0OjNC1QPHSWMkllgNdg6SL
E9A/PMA5HzbrzfFgfDK0RNe8p2gtQ3vOAM28B2YzDKdeqEJtwvWyX6j3jkYvU5pejsEikY5fwpn3
3F31I48j8dpN/nVrrha0bfufU8Er9ofoEoks86T8Y51mF8DrlAZjGMA2HmxiW9TCp5c3SollX33e
irOfU0orE1Vip2aaPlVTR7BF6DP91aSuNHfde7EKZmOgzmY+z2hL24Dz7QE2UBiX/B4d6KFC57oC
nMHMHHqfYx0hdJIhLmU+CTJm9QGAuq+rtHYvad9y+3qFxN71alPXkZg99olHLHarF0ZuVpWIBLcn
4BmfKn7z0QlW6J74jVOxjlJesMKcglgrhMXZNuZV/b3Uo2/58WOY4JofocDtRDZDOt5Kl6nLVl6x
XoK6+dCMHLBnH1MU8HGc6TSgaXS8q73osX0+3EHxnxzDJ6Qkcof1VY0GYGyTklqfpjV70l48XUvq
gDod4daFtdcqy7U9TPhYwaFI0MSdgwZNp+CnKSnrXOfAttqUeMi8gPPr+dk/W+opiYwFkw65rlVJ
TslbGlhvVRYhRWWtlyPsLGMQAK6ho0jn7QuKiEaDOnvTNz1b75o8806fkgG9EFLsTwKBCT22i2ys
zTNj8X7oA7ZVUD6EQqksLNGpXr0b4mNOjD01GTAu3Z28EYzQ7EivUwg9JM9J6SYj618LFld8E4Oi
YzGLy4Qkk3tnu26O1MxYHiM2c7eHYFTlV2Xs0L2q0TiIIWJqfl8ykii7njI5yuao7Dee/nrwtapH
oYTWf3/WyaKd3BAuEwwUpT/GJ1yAJbxuc5uwaIxtlYka+h6EXNigk80965Gwu4V2OhJR+E0et422
3zkryhe78D4znYfDThs/SdvejXuDSvajT22jzSpYjBpmGT9u325RADwDvGmm/8z4jrgHj+Y2svbl
EsPnIdtKHLA5ViblXqyH8hfjoJFupo9Wkrt5cfPeuqwyyr0GISzbAUHVC17A0ixv75ZDieUOFTDo
usCgvuMQCtodRHDmBNkkGb2CmryZ1zIufNMUuHb8q59n1NHN7hnDdfV2g5CI59qn9cBJhqSCaP8y
raUAZ9vD5DKymmoyfZ1QlYOn/VgJxjlVc6bGm3RpUa9USYUriwMxPfgyicGmHVKsFqSXNykCKyd5
Gid7s0PNmTm+bE/49FtYfMe4gOYhIChIXDoQAs1stBmPBa/iXBUSw7jUWRhEb89n4YfVCuFeOytt
QK79/Eq4d/JyKFNOhlvdE7CwttudoQzjK++ZT8wNXLOJpJadCGOIQ52bwUYuW+Fe/5OYjQk0Hxal
AHECSDzyiRhv0GAMBHFnLeLkbjK6GCstXQ2QfiU9L8Zo9NydujtuuoJ2NAsmUTOkuNjymtOv1bz4
GqAh+J4svNdVy8SyzskytMrolIpZEI9OMPOHfzvTWYGCiXhPNURWuHL2Hj6a4vj1LPInKVpGRLKD
/6VoHwl21NI0RRBshQW5fST63qr4QYAkpcNRkYIouvtQ9WStfNStCVDef7CQeY3N2uuiKVAyajQu
t3L55ic6+l1wq93cFg0kyZT2fQFEtjjy4cwf6lKfpiIomTjZYiOr3NV7U2ZdlCazJUA8bcXB+G+Z
pe0l1Y9piTrOLYpqpmJlq1qpbORQAPoBpATY+93q/DzUC/6JILgkomDIgMvunNQn+cd/7JHptgMo
cjYQ1NHWHTN0RaHGChboBc/BJ+qD3fWsTiMDr3cq0gCTupCNyjQdEwR8giT/MTa2X+8kl5soycHO
aYRojgUENO2mKxy0S6GbZ3KN2viOYHFegdruAGX3irEjhkDda13IhFiEOMubgM4sdnY4mrTZkCmG
ewy8lzl5Hz4DE1ODN7CKA8ebnR3tM86bhUWWNOfbmvUaRWJ8mi89ZXa5Z8iVzM7Enelbu41hF5BJ
sIOCG/2ffwdi1eW4vvLAZITMS7iaYmv+zW6kXTSQh/IGhN+GbiuS6WncE2sp0NYpyT9hqrVc9CLR
5I5dU5/ZAjfVYQCr3vCgsn9Y/PPeOVnZWnP9qYBtPMvP55c1ruDEvO0u6DdFLyTKjEj6qlp5B5lt
PpgyqRUTW/hH6R/ZvghMYsQeH6NHEMewtOEVaiKqxCCGuMR9kXsE79t1ke20SBqvuE8vxUc6y6yD
Fk9KeUyL3M9Va+8TpxqVS10nFHR/K+kSu7mLz7zR+iplFmwPaKkohrIKjLTpzYwigFIhkZsvTAid
YU+fJLtMk+RwskBIN5d3X+z/zeYIwPHQb0pSRuZ9jP3KnBXspXfUVREh7XdY5R5001zCqMNytZdc
2BDlISb7wS4ciq3T/AmQkcmqpp+S2AtetypW0NidkgS+9HIGYtHcu7TZFqNjsJIqf5zxaVkEqCJs
Kc2NW+CatmU2C0jULdqrkpju08A527X/ir5pTslRp/tMJKLFSU4wRRywHFP5D4wf5SYU7r4KsZti
w+fxuCOzWyUOLVEvZBxp5F2DYt1bZ5opkFWJMp3KnCV50Jqw4YGumkc8QwNcsG1fV9GfXyNwJNjF
RhLfRB0+BpIwHpOYNezLkq+2xnV9Rr/DV5RTnDbatqSxQy11eWLFTRN7R/lo3od8YSqI3AxP9gj6
Cs8l4g252ahfcSnQyJOwkX3orum2ZpxN0sjJGxrnHoK1DWSLFPHEEM+SfZsLohF1ZYD4zfwPHNgB
7tzHqzPzApY8XK55gk6+BBGLOcO9DxOFJYJHbUIutp83EYyBviREhkECdb7N+OeAGPr+HdJP2l++
4tVEhaB00ksW3AB84r//QXO36/oAnJ3DyufxDV29imtPU4ZDwFC4liJlaEEroi53l3+H+uzIYnJ5
N0y6qpZt3Ovpow63NyTLUoN3l8m5kurw32ds9aUvl4Ltq75MJfDRv5zf8tlyq/nTpjORVCRkBOLx
KKhYFWYMw2r1w14GsvQh8qL67QbZDKbWjf012MlhQBhPRxDEnNyZmO+HeGC6uR/UrMSIZe4cycPx
by3x5X79fbKeveiSqB2FIbL5cto3KxIvnN7oZrmZ3P8QxIE5xwJz8+/6CRfMBJk07A6N/OrTVxTV
lRyWA0NQqCZG7eubaWLAxdKzTx6l4zyblxdKEivEbp0/HgvIegZHvVJABMvILIkeO/59RPtuHsI0
BkEDo2RmJGTkfaaNj2FUsHHUtel9lmaclgVh9umLfEc0oNq8W4Unhj7fnAWuBESUcOQevWRR/rmp
fIO89NG+UFOFmTYI173Jd/AIeV9k8WIEOLoprqw8fX8EG+/s8yDe9yQZIJ/vZzGuoXkSvDMvGiS0
gRBbT+Yt0QyJqSP8/krc1oq7NdQ1sq8VjuXbkuSd0j0UOIZoDHxt2p7r6tAJqn4l1f38b/1gCphY
9tJ0WuUt+bPbKXoqIHhFNKl0AodZ3obHn4EetDzDVXYIT0r32obx/LrvAoEVdoMkIylos6TbZc6S
ZuwB7VdCN6ZbSBoAx/B61KcyTheq41j4todsGUf/NK4zVE0lL3WCeIjPwlnmDrhLMkxrQh+x5lEE
u3T0zj1P6kvkpArgVGktlxZhXFaVBQnXq8l0OPCXzGqpvYZrcHQSW4lXijdXYUqYfFJ9m29dvTR0
tmIpVfqRO1qykYUjidM0BndFAKH6/1mJ67due5vbDFfd7UW7sMnTHo3wVIhCI5qkusiU3EN5IqkO
BHAGsUlmXWhy8cqjlmgmhogTFULGhg0/XairiWyAiII2wfng+4XQztNgMozGlUr7/cCZ41NDAZIg
glOuasEUzltVCB0xqH6Aah8aN5cf/IIK7gBwHn8j8DMynlzhJvTgV0lrarhsR5zIBLcQFmxxO/Ei
7KGkpFjd8Q44jq8os4+j5x/6xM4v9DwOMlfzSBdHUd3jV0n84sg1fvZfZj8qdE0NVJVrbIKHQUZ5
shfpNXXpL0+cJRRa281oJPHJ4TOcM7Re3WGO7C1I6Ew4b+2BBrO2Ov3zYRaBvfFPDWg/eV+TTgo8
OqPmnDZhyNJVqJ5BCeFla7WJ1hpEBgwSesAhksi/wzETkLRTHAs2trB1yVuhlOAOb6u36EBmL7gN
18T3u8/MpH8aZ4ZSB/aF29pLrGZDtmJDlHvdHFpo7V41yjsezOt/w3QlJTeC6lv0Jz4qB6eDfMZ6
ESMv5ZayMDooXRCEPS1oCdTih6vkMRYIvDm4mimFtgLYv5fUxvUZtvJXCN4mwXrLoqZBSKfAmcul
Lkz+ED6KLrOP3qeHWDTdWiyQyBm3gGERkdnI94uwz24WT4MCVJOJ2e/fTzaAFzikQoCZoGhFR5uJ
lsyNrW0i1NywolKq7hpLNkmDrhhD1hg149nFRk6UiaTLPFCisqnJ2HKUFc6ndBiYKKonyeI1JwWR
86Mntj/bB39Suy56WSjjorB1FSTQXecPhB6ctalcuvgkPw56Htk4Ko24KN7DX1rGwGZlO1TcX01T
h29lCBhnTGNo6H9fGYf3BUV2Vzbq51AYyqpD+e/L+D5511hUtAc2FSDoklTBmTydbo9YyMgesNaV
DBbl+CWdmY3voUR2NDpaUvL7ieCA0EqNZJNrcCDbMrxf4oCGPtmIW50XzZcb+73LIbu1AmPxpdY+
Pb8vOtpWWrnokZghKhAUjLMtjSdzTsbxJDT4es47/PFYl8bMhgMnju4hn8BIjJw3rew+jZZaEPUV
SqsP2K0swlX0pyVg5xy4R2uTaJUl3izehsZpZB0D2wYVjzsqj2DYU/gzlw3vw2CuhOK89CzMILeo
z+CgdK999bz4ztXTqvZTN/Oh+1OUdsJ79kGjM0WljIaVTZ323f6uNLnhVfLTFyPMpP50kCZu6nYM
TLLA9dq0sJDg90XrFJhcjZIRsg+plU95aTPQMuNvrqp79WwaphUKPwgFSFLBb9pt5tZkCvwxclJx
erfhc6H/zp5Owh6208BhjePpTemf6wN2bgTOtHSP/FcYxa/Gj8lEo3XSvR835m/RaEbzvZG2vxBO
lkyKIGEEhdV8UVQYqhVd4pyX+2JLYrYUH+Ex3Mca+AW1bR7bcgBn3dIBOTOsmyRWhDmyLhW14j4S
8jWRpi8SKScPEqBZ6Os4vyIyH/7EIzeYvJm0fkvTxN45QHQCv5TJu28qHGQfD2Tk8xNXhU/bh1oe
Is6QHc/79+nejR9HfNj8hS00riSnQW2Rgu0vgl8GjOE4NtPMBtg7IOPa3t3H2RuNczSmWfInM2bh
geeGUNjJrt7JERmCSzklczG1aS8bF0PDUfRrU52B2rwzRl/pCo3cW3glXHpXBnTVkUfeE8fRxJ9K
FVLgMhDLVq8hTLM4r6w/+KWm9phqR6ce1h1PMY1p+Vlu3NlWw8AeHgWC4xg1nDPV6EORMSmtwsnN
GleeO398xS5BnIVZoUu3dW/9NPcrrFEZfifNkZBTH3oAtImEVqWj8+pgdys89u4XOcqiwRkykX8v
xPOfP61l2Ev+cjjkLV7Oof9r0rmJow8StN4yikZRNB24gtDqNqB0vohgu20TeAo0R60DFxdb5EoA
O01W6bRzCRr7R7Ff7ScfMLyUy7CyNggTIBcZfhtzhmXY6DSRBNoXGEwat4b/knvfWrXIHc+BNsYQ
+5eeDsOAvseOt5vLnKRCvgwzkjs9/f8tKQ51vIXKTqdtsvhmBPZy7v+i+SVfiA4g96yGEMDiXP/j
jY/QCVQ+MLwEbIruZWN/ItwozqnRcOjLKi8Zoo/wk/iI2XGZexGxsFMuFVOcNI4sGt3OvRgM6r86
k/J6uOjHWrmQzsapT0fthIUxs5MetV96TVAWYZ70JmFCdfwv2vOy7DbpHRGEA6Tq8MhYQAqYrmDY
OANpy1yNJqujVEWp/fUYvkiYRMRtKjNsMK+rW8l2WHphA69VPjb8hrTMsR1i37k2pOcnVAxh10qh
d44iLyX30ZVTo7siKD2n3JznFrHsiy85sL0sgKchkDP2a3CZfVh8yBToGL2vA2Dhaj243ZQAbWra
SQo+J+kMo9uP2B/xU3wFZq2Mi+B1Lt65si7J0nWbJ/4OIMA9tMb4ztxIWOKjPl0EChVTjNoYxZ55
1mr+LOvGWxWr7uyFtn47SDL1s6Yvjp3ihy6FilHeKspBYl7p2Bm1LIa/MQAEvd+uRToaoALcUdSH
BHOWWrPxp6Bi7GGHX9Bzey62gEzKYQgiFmGUIGTblWl1gMJDE6yBf67R1YCl0epgoZuOTUoidVgP
LoS2Zfxc5s3Zpnn2rvLaWRgw/PuSC0uLsrEdwwznMXEPUxLI3DjpGy27hgY+iZs7lJNuIIf67sBF
k1o8V/d55UGiu6Qu5LNi2FEyYBNQCsrO2NvQTQGX3kK8xYGCUDjoyLf3q/nltC4fOQoqjrB2ZlDw
AcRDh/k+9PqrUaBRAt7SPRHPTT/3EvuEm9roAGvkbakgWV4sSwsvorCjGN5Lk6VjDZKiim5AybN2
n6wV6K5dwxj4CsEZoo4MpdXUxZECJqcpr1i3MC156LE9HUAaPQnL29x5JpJKSB0D+k01pE8Yv2De
Ba8YXFnAqujWYecfLnOgJBP4ozSECmQB+9L4Ks7qoR9rh4EzfyoY/rop2h0QQaVNtsN7A/iU1soi
iYCak3zvrF4s9aydAsxK3b0nbXLRtK0mDuQ6OFQkQCvuSyQiScUfH4TevVaYqvYo8na1WNPSLyLk
+uhLO4XZlQEWgpnqn+rsbySnbq51cmcivchvRZnA9y+kF8S+asGRxq4Kncu3MaW5tQeU7cixGN4o
72co+8++4L0T3umo3MhT2rCgUonU9nMiXnLZ/CzGVtmyBL6IS1ySFp5JSEHn3I6GBsLe/8Ek6lzI
sXXSJWwlzr9sVUiXwvlOhXSE5OZaCWSMiiyVEC7uSrCWA32Fo7Xb+UbpDqy1XVg+R8hwTtKuHx5+
oyacmG29rUkdmrb/loyJO0G63X3DghemiwDhzOzcjByR/8m+1YdTClnREgsMJyvLW3qHIfm7fdKS
/NEOzDquuQ0HO62PDjlM5abHtoiaCcuREG88jwcj+P6T0sil5FU0UWSu7WRJEbIcf16fTQJtSQdi
mndGaVQJbPpYVqXzO0og59rEX2HvbyRBVEkIGRUoOxQrADKqwDW1cSH5tUNpB6fycCI8tHWJG3Ka
VnQtEcze7Kj0CtsMscG/T8rTTsqG3VYiR5oVPFfYDc2gHgY9ahNmoBFRV2MHQp+GgjmxuX/vfKoA
y9PVABsCy3OAxMjhR+lMhwIb3hUh+XrugWc7vWxkBlV9IqUWZTj1/SvYAdIIvWU8SlrLIOnEEMte
Kq0y7K57j/9DnV0E4cOoVwe73UppVJ1OpAYGbwpqwJyTdR7I6v2FlkhQOptgm5pYSeYjk8is3GID
zWLGhxQjaqmIMLlGmY5tJgP4nfEDnaSNKA7E+p9+JIaK+KmSVTl/pR092NFSWEVwBY7liIi836HN
U64X58ouUKjzGKZr48+s6/sVCmMtyJf7jmha+wPftFMHipiXiSvnhbEX7fjfv64pg4OJerkctCYi
irTWw2aT39We01wRwfZEGYyK9IuDw06jNIeddzsP+TLMGIc312PVUfKhxbi2GUXTev46qlpAw39J
o5RYmamY/J3ae4fqNF6kryxTpYKguYAz4NTKXygxEE9R48SCoEQrXQBs1Q8r5p18o6hPZ4nGSRNc
eoiYMmZD3XVQUrznEi33D2H5QwNeurT5j7TwCu9jLfcE/k64XsgQ3TEHPdjclIdnMCD0GxZxJ2ho
WQybqccjSCfZl+cvrSci8E5NHrWRfNT2uOdkwa/nHimIWUWlJSGOvLaWKwqYMYMSxglUyr3pgLzs
GmE+gLT9RQFPtWeXLKgBmORkBZgcXtj+fSC5KlBovOhNS95+ZgIPWyfJgddfc/nF4X/buVMqUUA5
aU8QwF6geTyc+yjDD4ZLm6aPyBkh1N6HxUEDA8ol+rrslcZUibTMxbjYbnjhbBsXnIjdi+o99G33
hPBvw3yU4TLZGB+IcHrE3Hh7KcA2QKKjGKEx2iI05MzbQBGzhbqUwIcBzCNdJIoqTwUADjiR33nc
SZ/IZamiAjG0CcGnS40NgNRt1N9r9k0d2a4eRn70IZbrEnr3NgLIJueP0Yt82ZcLCLFn2XgtWP0E
QDz6SkwVDrDhVbfZdLaBMcNmEtICJ8veE3uhdVzjDymh9pKZJmGE5W93SlMCxkJxYNB7NRGeMpVe
d9xAsqvMpt289n2CCwfJOA6cIl2Q16FSXjdJG35rnFLuxQpWOr8gCy9HciXy6w8tZk4KNnAbYvf+
WLl4k89anH6QzucoQkdcny+38yNeaq15BLS9tSGzgYpY8P3brr62ymzRN7WZ86dadZPtWcnLsqFz
uYsRa4If1Ls04z0N4xxcUWgSTi70lNsh6nsTwR5kT2odWS1D0GoK2GgvSbJ3GdQhorHkBvJeyZC7
R8ooBl0oeE2y7jgbXl2JhUzr0TDtwPjNTJKrcYChXUEkWmozncjgRL2V+vZfI89ue25/AKCqvjK4
jLHvouUZnZem8NhD9/9DAbbUpXnMyJkz5qqDK91CqCBg07HN2ABypryBnR1DrsVf+IPx4uEczXr/
yl/BZRNJLYej68PS2THCQ45o2hetzVOcPlpk2E5Iq7uioU0RAwHRNw6/jHETiBrndQK/s5ruHcB8
x3BkA4YArCEVBTfDQEkrUmvo546SditQgaCMtlDMjGMjrk51f7Aqcfb49l8oy9byXd9V8ZNqa+j4
y/s4QLhB9gjWpJtNFhsdcZJP4YE38SYJQdSnSRBdk+QrgkX/f5Y5Sl67MPvmgOovQmVU3MK2RZfS
qXdtHBd9wwg854oFM4NOmPGfQ+sbvJwS1x5olpeW0Wk7RpiLge+mv+1HL11Q6mpkuKbnTDDQtaEd
A8QjKE+M7qtMvi5w/coUaVw2BD4fdGdwfK9gD5A+Lop2R3GAiuJMX1zBdgkJfYuUo80iwVY4k6Fu
ARsqoOKmUwsmCJMAU3MBL09OieMo5XJ/LkqyQIJnHX5ueiAdC8aaYLwluQvGNtXWlT3XD+qb6FKe
oIK619BHC36fkuB094scFffrjJ8gQO96j024O1qnKngXXDoJJyPkD1FoVofmyBlrb4NMjh1+9ASw
70qZHHBwda8HQ4CBCQnNqeXqfg+eD+O2C4d7JdoFK7YH138JXggqVt92/Tb6XEo80Bf9+XBHeXwQ
miuXpu6uiNUUI+w+oLai33dB2NVN3V1xxuNwkNySbnhnB0CzqUhe777Z3P08iYOLUE6kfVFgLJCY
rL0fw7lMBPO3XhaOjtA/7VdYPM/1+qqDV9jRDLBGT1Wyq6tEAxRePfu0hZl9PmUOGLHscKB6mP6r
6Xxs0Q6+eFfaDDNIxlFeNmwX4VsB3hnP0L/8GP6Z+wkOGU8spkiDRxQWlAPbp+iVHKfApSMwg5q9
a0LqoXzVxzm1YviJxCVBL5EgiolFlxv/ClQUEgOiTvaW7/7VxBGmxSVjH7UrJMp+iMslaeC87u+Q
7+LcC/byppGRO6p+/TxAklvHjHSwajW7BPoToa5Az30V+KiLk6jDT+pl/Yx9clcxsgoYGt46UvCd
ZFJ+SWTB7QXd2coaJGypJ6Vlfw4c30xIBmRfAL4/1Bsa+xmHdlNYWc9WS2WxDHDMSQo8uMEwDGPX
5G97K9CrAjSiF/sW+aBLznQ9DxcWNGfJW8QwH8CZocb3pF4ykDE5ctYi2ekx/9kZ2tJrO33zfVsl
zVqEMsjAQqWD1eOE0d2FVf/MpduPIPBkGJeEUnYbvSsPqIm4AsLVoU2Hw60Gd+AGZGCkywwTQtNP
BUroQ/48eQo/hMuFKWVnkE9z7b5hAjQDsWW30MANGN4OQv186oHalxHvu9m2bR8vnSqEVKtbpwHB
+a0/jao8G7q2wutaW/oWhCsPSbMqmvCo6JZmc1ZoIXicpNyjd8LR+yu2rAn4gKxrqtfVFSjs1xIp
PnC281Tr1/lp97H0aRC6Ok/CuB38IIL7Ad8dunHnQ9z/ba6mwy+fKr7FPU2r4IXJL/8AIelcvLmG
n2fqvmr9L2qTvsultbpoAW4n4gHQiUAoNMxEtTOOpCb2gaz4dZMfeR2AZWm3PACsXIxUk7bYEgKj
5oqp4rLv/jeSO4+HloPIQAd35M1N792/LyN2pxzQRcNlL2DmbzP7p7pFy/bbk79DMvspFwxgXNMe
M7cuQ7acOxFBwmytQDlm9Xd6y04lwxxKtgPcg6WHKjVj0jpfCUkTUxYSVdPUZ5rZdDq8318P3oF8
yD4qOHdD4AOS7nU/ROhZ8ZMvSBSK2aHuySpH/OyGLjZx+5YJUAaItU07T9aAk+wVO92aYISMq1PD
zO09Sp/TFJ4CQN4WVPivqTN7yqRT7uQQ7UIll5gAyy1FONC/K5OluXqGsjB63GYE6neKx6X4qTql
GsUfraW9n9TJPXPGwYK29WeI0uH/R2E7XVX58B0cK6vu3I8hxBW03I0rCVtZW/8ildAvinzy+EI3
yxJF9DMjD37w1y4VpSkZWrFx4mYGSlcC2cMYfGdgSWdGKBA6udloTQpIhJHjIBfYq2J+Js6zEw4X
f46hyytDVt1Xji+9EYuMq/T9++MbYlLKN0uwC/nzKIpgs3lMhq4nEKZ0gVfm/T+XFVEc9Zlyh+EA
Am6hUVDq/42TlcqLd3/xxn1L0UcrWsmEMKg434CgJeQEd72B0pX04R/j7FQ3D7qjCrTXvsAmvKUu
6ud/ECetPo+gIPdwiiGeaPQDac7ekEZv9EpMKNnRdNgEaquLQoVCSMB3iCX+Wez0vjuNf/YIKeki
op3qbF3gwP91QRKpzhIUU1Br785K6i79rdTMLZr4JIdh7NuHVckR5X6TjQ8bC+p4hBm1g7EyDc5d
n+JGJ7/gaBTIheD/yDwb3S/Y4hLdrEUeVQD4WwDGS3/0JEcvgGX9g+Fy7y9owUSE3khuI3SVdoN2
BlEuTisFsBs9zV96YqohSURrA8ROuODVKCyi37TF8mya+UTw4TNIPCYAvMqp74y47IYUudDfJJKs
ILr/Q7RR7YfVDrY7j9iqBoRzXnauMVkBV9Oyx2/awpQ+fUEbLPI4D8NVG0S4yfRDvxA63h6gx2ku
BN9cyvX6hpYSkHmZKt2ZV8JfeMr0DgugOai2oXSh7lO/oIRagFY4tiTbm8VwC9oOQdQhtdpMO3x1
U82pkeW+GjeUOgwI0u7VZuC7+1I98hJHWdiAFkDaMvDZbFM/+gqfA2spkN5+k+F5+D8gdxiU9sBs
aJDT63eY0daeWwKQPUv1T9ZoUXIdkPwGDe9onAGX8CtWsX0ubkreNAfAY4FVHTU/koSFE5mwPWRg
YFNKy9YbtwpgMoU8WUmW5v6sDVcoKBFFFRkrYj/S+7pIGaw/p2aaf7n2QvVw6X1DJGugWyeeh4O1
C7NC9XUoniginiL/pkscaQWlXPt5whLBKgATQAQeYFCyzk7GVe16uqElYkRxT3q5P+cKKmc9EpsS
yKuooMfT6T3155/uApZ2sTduxCE0dE/ZQHMa5DoACnNFhyXgAJ7UEbfBeY4WMV6WULByuFT3tYqQ
TfReJprEgZcATdWHWfd05ExGFbKPWa5zy1uwlaAVnxPwX4fE1igL4PLv7A2QiT46UP7EVMhYPgdA
fXMhOg6HSNdNv0dHV6QqMisXyC1x43GIKut7kp3ymkD5b2MOQfi33ltmoHAj858zZLyRa7FkRsHh
GcryZpfC9jqWL0YE+11RNBHTAEbE/hl1aIcA1qm8IoeROXCTMJmBrIV9pQaFS98vSt/oQlfwTWV3
+/IeeVRRHzMhtxLwzfBxql5w5hyP+pHYv9SFsA9gJtCWUKmR4pYYJJoDIuSv06lfv86FUlSR1HP8
iFqW+HmZEs3sE3pjsCKMuWOqkE4mfLhxFkEAx9XzXiqDedE07nvPK48jCv1VgZZp3uGFZgzr75SA
+svXqxo7c0THGXwdjJo9ilyCzDbai6ywoCa0utl7lEHS2aVYgmsrJXYdOSSqHLGr7HgaL+H8XZxZ
KEXqyax9fCFR/hk7DnV4HOV85ykPZDZid3bac07037WbVFvZJQKIOlP/KeGMaUs45ImmjTBqmCTo
onT8nmu6hHRp3y0LGd1wKYtYkWKkd9h9dAMKYo2bb3xPmZE1ZqwOce9TJxIv4id/NDiPBhi/07dD
RTc5zsWvA72xZ/dKYN0yIQDd0eLChzeA0qYdaB/I0zOxe3qulJEnkWCVrqIMIKgvvTuXf4vha+6k
LfFNgfyaPxWEfMMcsuHsmdzl1764+cGyKZbRpsYPvgcn5WPmfSbNk185HFwK4fXkYGNW43Oz98ZD
P3+jCRMOv8hoswfll2Mui+Of26qv6Nxqh9an45YcEeMPZSzAL4TAUWxHfmksB96TGBJmp5qcruAK
e7NLwCrGpKiC6Raonq/mGrDI3Zn8ykhvaW8zR7AznSWez5e05HD8tTdeUJCqYQTB30+9gYG2aP90
/Hdlapm2fBmRA1L2+/xJWqPlin5L+a8Z8GJ/uXohM6JypkyEF6xfAPNHPu+dfbPB+dGm1TZQRlyZ
lQHUP/+LgCB9da7exaGsZ2EqJkoCudI4HGXeaB3TpXp5VRPYjrYESbDSGwjvmg9tk3lLdqRkkYjS
FZwVWL6Ay+HBiRDeMI53id4JlCP/fVji3vAjyJOkBEP0knBCr9G5lLT7b1sZPVLMlGTf9c0VZJyF
9osZoB1m7/Q1hRuUYSUD4ry4H+mM/zagQZcjA9pL9o37hcZL6i1kbeVyKCMLx6dCMyz0MaOXFwEN
9Jpyl6TXzooCTPda1De75mk94AyqBbBTCCj//lnIT7ju5Ra5vS5qssxtBw7VQcFXtH4/9m+PxT+l
NmIVfbkXMPXjnD2NQhthICjVmMQRplEEtZJMJhpIJ/YsNXtj0ANUoDeYIDS8+A96azlO53K6G7ef
plBJTfiDSG/4dzaaMOohIN6Na5LRwvHhGfIZijDNgIAZKbaAha6GSWWjnwy/J/9cAv6oqgI0JYCp
/P9p2QHkRsTiTd9tKkHiHToKGN9HmI5TUN6sXUP593Kvt8qPhZk5ENXzID03+n2F2hA9ziCZBG5U
l9JpcQDE5vVrpW7+9esMjmxbsThEwrX+sLcYceJr2J7DQcXLoawvpUpPRKNsBzWoRRgOfCcgVAha
khrCSFWEmGB5xANV+saNTCkxm1mH8tCu+ipyiF3RBwgLrLREoTV6v5o+zKkI28F3GrfGsu2UxPyt
b+TAn619P22e8dgU/POvUZnqXV7Pzd31T/a05T1rwJVEGqJtAwlqyvTV8eMvSQH2DUQrdca0aH8a
bijNgO/m/LUR9KIlLSXLYsN8yR7y8lVpm69LFY7EMNbKUryamKkikMQE3hLJl9hsj6LDcqsT3IAJ
UFWnE4eMvjA0xSRULuyePdQw2EjJpW1KnaYAIizsRKexM62+ZYk6Cied9sYE7EflGfKh85hiVilW
1lVf85XJzOm+CZJmZx+3W73aLqqPrtyfQgJUYPESJ+eNCOkLJDfSoyZZ1BBlEpceSUMyy/STacu2
h/OrCo+4EpbaHak75anHPlLf2Z4nDEE3cwNvCb1YCXSlNxRnRfWawI5a2IGWzt65JJEmi1FIhAum
8lYkxFMY9SCAQnO8N+RoXqYA8nLl0Zd0YNTXwsqZ6L2lZZgH512RzVMZMEs5pxlEdChjDt++rrnm
GLnXA/hqS9eWJ5+jFKNQzFuLWYxIUaXCZogP8dxXTcf5fO12JYyZRe6JOwedXg5CCDnEm9dEgu2J
RTUA4bneq9yhAWdSN2wiLCOEXCuj6/0KwSgWi7zLX5ugOs8OgOar6tGug1dBGweuOtiC7gqYOHDJ
EdBYRU30ySF/VpSRrFGwxCJVm+12sQ8dFvgoOKSh2IrqwZ3bSkD5DUKi+qS2fDs83hpMX5+4qW2A
GXo9rI6pO7Su2redlwahycr59olsWLuunBFzYg42I1QDC+PuE6DhwrWHLKEW/fm7fhApLREoOnWj
klE/mbPdQmEc7QSPpn2fuvJARwBx/tsSp1raEAz6efwoA3nB/0HthDsmJ1xQeeKN3B7HEkfTdIxl
oqiG7WIsWa+3cxkvWswoDa/Z5a+HQiVIT57NhS/xNQ35woFLFpkJ/EtTzYj7msta+wRnRdarqpSy
Ibh7St3wIxqzksNwzbUXIZBiBWHsuxk+UaA+1bTxQ8qum1faZVWSdbHK92aB+/+2ozvM3PRzzspz
qO4wBxhg9GPH7Wa/gsoS3dZjnpZUOu/PahBn8AmhpoNhO11QpWHuSxk8uefR0ESbqUIC9dg42QSJ
zICf+6hHgA3xKLmyC8DGjxt/+FQjHtsNvG0xCHOw+9ulGU4GhahSvhDSe37Ey2d0E8OiO5cIy8Zj
1e1zcZ8nx2ON9IUzMfUL4bMeURrmOSnTZojdrROI0A+f+fVh1xRGjVl9wTkfsmquomV/OrY7EVZk
tmxfRZ13QRBwDmbzd7jH5f7eEYWRCyex2cVumd06vpsSAKNaW4wdRuj46swg6BLl5LofikTc99KC
kT6KAFaYijIyD3ox3AUynAZQeoBFYzsDtOyM0pdZWzrzhCwVcJskVIrLkPA+FRqCr70XrHp3KV26
bujhcZpJpWIND6mELC0uMh46BCPAMEDnpe2jCfqzqT0KRz4oaaAhyZv4EdztieSDIgaxJglR+3IR
Y1OR82kojqsV41aS7mX6VBNewCLiKh5ATzMh0bgt28U1FUFvgKmYnOUPxJO7iSFx4KMRXfsEOy53
j/EhzWv153js2uUR+nb5s4PNhBCR1UBLqOUfXsVphl5RODBaJnRbfXzCg8H/SQBWb3QgwbhxKwl0
J+Nl+jAkWnD+WUi/tLAdQMGMz0qeMMWXqBbmR92QlIDfWaxeiFJkMhqwrnb/Br9KCt0pz/v51UWd
bsJqvzR/Cqcr3IQHvt+cAnLEQlLd8XErjgSjB8yOb6ajddChX0/8T1iIh1xW9xQB77XrVMbJlHBC
mYlOBhcACpxpmBRAf8RBKDSWaa7apGAazdhTGuBt7Oiw34NYxRY99X6KSeBzabHlw953uscPDJeA
MKJzCdne8oRS86Nmi1ft+EZJwy3iPkPepW5Jk+ASlitqCkqrqbGf2IG0e+CRjRSEXAsxlT2u6I4q
NrnV8nXaueY9D4m8WjXkNM3TOPojtJKT8hb8Hpo1llvecbQY8OZv+1A13SRMF/IbnVZgETBxS4z+
lYjrGtB+XdBOjhLNBO2Z7qGpac+qRHVD0YzPBwLfLJqj4gAP+9e9pl2uh5+EYpGxSxc/gK28EmRz
ZSFllyJ0GOOi5KXFFmtgZF/jdzTJuc7fDD0lgM39cnBlBd4amWpkIaTuIu4CdXJzVk71ZQANY3Ie
g7SfRWeGmcrPamdJtppi0ejUFl3aWSLdfv9/Dn5MFuaTwmsO/ipDYBf+ZIbYr2ET1E9aoC/MUE4+
X3LDiAIw3kYKqY2tDCaEkoDfsjC7dnTIFAe15D0+OZVOm1oJOUM2+uOw54QtMRthp1vR2ftUmPDR
wVqbSGM5HSKkkhqHST8rzgxN+Pzfp3L5ZQcvvuJz7US0KFNV3U3Tx05h2OM4P/rnz/bhvf1ChFf+
oXi31k80Pu/ZgUPxCx4J1BtT4ouWSf8HQK14h98NHjbZkZnb/q7zdxxrluAu92Fb/cI9J3rIyp3c
Gl/vaDJUS6RiwSHQi86ZYtUTFZFSHyF1aKULO58BmrlvSdj2+rOy1gBfJAKWn+DInV2e9nEg9gRt
ozPeiMyEQ6pBiEBf8SseKROIz3oUMIfspLfilKCU6VUxSHLHrSgCgfhQeMlPwzAP2sDSyudqSzx1
OYncQhTqUDFDE/MciZiQlj9kb6ZsNqQ0mfvdKI/WYbJh5nbppH/PhF2lwxHCiYQBmpjN1aw47UOr
p68bX5Kkyo3ShyXp9/Q4tyFmZL/w4/BQYwI0S1iBEIfNJCku3Z35OzeUeIyYiYRia7ndugLnxk5r
F5wHUVofiHUQLLhvoXJgbrb9AbmpCxJE3FjKrjYppcggeFwQ+49IXi3p2WEdTWwiRtYrzUl+eaFb
06LqoD9YvOv1cVDZ8RJh+G3TZ7rcZbZE2cwD5nEErOXvzPI4CdsOuhe1BLU2ygn/1D+Rkp3T+2CY
Y3zY+ZjRSoFBL+AEm8PZFrFEJEkdpgxS9dQHdFbHO0yXE+6c5aYutU9DRLXITvMYSzW1KIsMfRor
jLwK9QDWI6ln+DVKXA2ORNrTScKkXA8GBAGoE8ZxZSibNlzwTQ8rCkd1qL4XhTlDgBgE+aIs9eQ7
pvRR07e0Q27igL/m/A9QkXfswoDR82V/vddXIXq0jhoMioDZwvadBcIAwJojbWXy+RGgkq6b0Nl0
UWnKnCtbpkmQv+bzSfPY4Z7Q3WzVQZYvKi81idcOvoRjXxh4AgptOu3z9W9AYDJfwWHqo4ZfrpDe
cfMFvJQSRUMaSOFCG6tEBiiLDHGODSi7cAhcfSU7ODtuDH7Yqyu/STsoinEdNzEuoIemrFmp349J
hT3jJUZsnszZLQ621Bo7Ntr2n3VLbEZDfhmPQtJXqsnYI4wSQ+rgkv89aQJWH2XuuZ7UqYA5/MKO
Rw3FGjj1SRslhwhzGz/5tEl5XghZeTLbW0iq6TfONEJqjodcpooaJrw+i/uKl+2ECH5ekvHvssmH
MbvOcfHnVv48FNzreiVJ63az0ILK0Rbw0TZsU5X2wjj1GXBVRBkHxTrF2IA60JzM/Unp7tFhjP8P
KbZdF1Q3bWiFDysWsamHbw7HMJJGHcFxsblc4iHGKTSllfjFRzAl1n+yTP0VYxjaqLKTnviUAZGU
WYCWDnucUwolr6RxYyw3bKnH/S0LajDhtouOa7kvTQ6joRk+JslamCP4+mlpFE8MXA71QeIzt9db
5Ic5yPcsBHH+8sFeKoZBKjagGGIgZC8L4V27nNS3JaNRsgiXhBAls9figzOR0kVaStwPNgi5SO8k
Wpo654WTwxcvHt/nZ9h8tLpU98wPs86qvQ5eueU0XQfkTPpi8m5nAO0RnnNXroJ9nShVhqSJda3P
I7MIls5NYqvwCj+ySGyJvnNoi137r9LwvFoSCWIEItZHA4RbsIKtTGZ9YNa6ES5SIiN3cmIyvs4f
iOS0QItPtMYU2+ECjxAWo44TbyRHvpAgqeWpt2lkq/EU6FUD87YPxbV1Ul6UnWxaF5lpsf6lT7Jw
uF2c/kZ40BN2KcJtmyanroyGZbmCT+8YvpFBSrkiM3Is2XyD8jtw4EDvbufPBQ0frUDbM8+Xe1U9
MsF8HytchnBqJSs0C91gzxOB5to3Kf9ITmGUfsQhcG7LmSIJrHTJStEbtUpPd6aTy2CuLPlLezZ5
4rIRqA/SM5suAdn6/sD8ddl0HtM42W0hMR0raSQS2yOM8HxDgsuApwgtyNI2CdAjZfmuwUU+ui+u
3906k2YD6XBmzSfl20E6YKZOw06oEQY+jB61xSokp6EIAkY/hgUALYklU1ykAgY28BX4waNxlOEs
fjWp2iPMdqQ6oJ5oqcC5pO7qpQq+Z/hUrfomJEtbvTSARdOo6UDlmC1s7JVXTesEWxmHsLUK6xtA
6zC5te0YYW77/uEq+3jGHE2CbEpZmomX0gdf9nxu/6gWKIoxBmIXrojUcX/WarKJhV5BlwaHxejj
+4/RkOyEKetNRPfu2CfejEosphm/gCXaG6y3mnYv2V1MtqRBCh8ilohr41AsPLwh7gz79s6QH0lb
6Ci9zC/un4P+RQducn1ipjoNb49OBwTas4/W7f/ah/I+WyebO4oCCXp1U8eGxpijED2G6l3UbhN2
+fVwN9VXqVn842gN0Etkb02hPOY57JXUxXdwSeXJ00x98U/wxwNyl8zR/DN7+oRb3g7CHnOzlenY
Kx+7o1/+61Nrn6vkH4ts/9O4oIe8CBks2hTvNUqHqVwk9/Og0ZwOE/nfzquomHm6nVX9k4Hk/Awg
F4BUZEVZqGn8ReaHELcQM6lPB8699q9+3r0r6qYgK3JKahwDAtbrUOBloutXsBTuX8aOy6/b6aCS
OZBpeops6k7VNLJqyT3rtx3jkcWnSVkye/WJVUuaJsqPZ+xumnLdCkj2tzGMXC/sRAmaScDjqRNQ
0zCiv5J0eHXFLgiSSkCmjUY3O6Yo8BtkmuDsDRXpwHgSuaWQt9uvT5fzg4KjHatj2Rz4HDqg7Bgw
w3he7cfAubt+h+Ik8IYhFPYyaLUKVk2u2tQJz/dFaJgigcTFIMvBSZXhMgWyVZS99gD2loqlAqND
lg6pwwxfoVJFS0K935syU7ktgFbvYQZbQT3kSQouQPPKMON+N0jUe7KVYlOjgXKhwAd3NJGSWDIZ
Uj194CDCOMemKjq6MvuJVrggPDaGgF5vwrU4yFAMdN3auxSQBAi7F9Uqm6qULuFSLXZkUOzty4LX
pfVckOZS4HWIuOV24Gtz5Q5TqPjNMYFRu+Cuh7zSijUhHGLky21QSIBdnEAL9T7zwo16aGApD9hX
e+opyO3qkWZRD6Db8FkseqozKYRJQz28mZCesU+vd+XFRNQXAQu6+1F/n4IlblrhpMOUsXfhvc8t
N+XME2Cm9/vlh6CdmZ3+oV7W1tWZ7cflgYxG0oJ7kFlcTQorcOim1UzAXNnUSgeiX1XYqeP2kWEs
JjtDA55n3iI26TkXCmR42CJde3zp69g6vwXPA6Y952N/fBVfdCSnEx19n+pL1zUPBM7E1ICt2wcu
fYQp8bZxujyywGGAVMqO0BqnXEI/APkQ+zx77W+VHWiIhxkGVsIYugBfU+CTqb8LRL+/zujdsh0c
yrnV9bBQS5AyYTp/sRwbGgMd8ch7KRCLVYB2iDdaF59/wy/SlYf9btKN4TrqrICpE2XzccnXK/Zf
xN1bH+i3r6C/t3k4AiUVFy2RMt909Y8mMTyrnU8+6KwM8eBzomzzaYyn9UANVNgn1kYSu5GbfJX2
7CAf+tkYSUp3qE9nrQ/Oml0VhkUcd/q1IWbo5Fnge0VJh4UKrXFQtb7TEdSZdKlWPwL7F36nHnjx
oyhlCJ1JkF5AgfoNogkf5BOgivLlXA1EAyRVzumvZRFd54RL0AMKPeFqzkqfKLE/9Roq/HbgQ59c
udBPR/1QBTin1sAxwPaAc330pc0WcYggi0oxpuvzi0vFzy4bnWoxQMAsf+T+3UD9PrPzqvyww37C
tE0OYaxwSDoIzuhOJv4jmKuFrajWp6ePVQ0Hgo9wMVmVqo2YIyGRCtt0CPvaa5F0rx52Ii75BxTo
apMI14fVs4UDdglB9jb/a7dBePSB54TSO610b9J6r2N0S+Ni2Y37E1j2YlOt8W5aXLO2IV7l+5pi
bAHxcR7+td+XCOC50DLMp64mHKLFLaVzghIJIUEnMvSTpwJOrcCEbHFhq5w1FulMrTRWiLNacRIe
Szh4ma5+OxqUxcbxSvuLC0W2sRBvio0W7kRf5XDZ32HYGNgmZGMMIdtRHfmqW8X8F8VXIyn3oBtm
XgY3jfSgEiXGGBafbHxLjGJZWZhMKHTFwSN6+0XCR95+7i4w//XK3drr0MVQ7eCCwcNyfADtI2hT
MsKZ3t4kmn3T1TaomUF5hcpCCAEbAS1yo37VcxtQfU+VIR7gEg2ZvUkz8xwVQZMt6iBTeztOvG+q
6DSZfVynDlN53fEfYmGeTh3DR6tZXRAs9KV2sYJPkk6aL6LUoxW1YEht+zxyigg1bQ2VX+wxlNTA
N9Fc376rJANKDUN47VxGck6kC7GGc2d3bPNhulxVvSuXu7xUvL1IKdWhLghbMT9QtTsEZqhSaZfq
N4sikBETxeBQe7nGhkq+3RapBRwzMd3odzFz+RSoevYL2+50q9YwySVhPXCZzFNSGthUiHoPc7Au
63IfRj3Tu3xD2jX6XhpMTaHD28a3Sft1k64a1oihScoG26dk6wymt3sl8bN9JlWVEq4kygKEOFha
tY3mx1+jcYonNV96ZV6BMfqdfTccZxOEY3BEtE/4xql6UKzi/lW268UTFhEFFeprSHclunqFZRUA
FVF7tCTDAzNbPqTl9ho9xDGz1gWsPBQLwpEfaxaFs3ZDsdrZpMpofM7IWyOSujt1w1Dmd4w+Dah3
x0HMwE9z43jZhMEbdSO+wGYqfZNmvxB604KmbvpDv9GtHOtnxC/FQyf8L/3tu2iF9HqHCflkpwws
Wj6gUmJTLZfiTLgX7SZzZfs/pJdUpFN8elBwVjOvzEdA6J9hQJ08aUgteMINWodCEudMBQR40Yvk
HHmeufE32EWKgWIhBvF6cL+NgknO3K+QlZmu1Jwdyc/vAGd1VgznM8T+2O6BVU0GHFj/5tFx9LAd
9NWbFOmYnX51doVHUtKb/ZMt9n+jeyGdTPwWe2JN03zWj5qexVoTktEUraz3kDA9obUveOqcpSEr
Jw1Ak1h1cX9N+ezkgSaKNqouCcB3XDiDYLtaPttOyj4O1Hvft0+/lKJDaNnHSB3FCaIAKAO2RjRm
lm+LDcO5PFn68AoxB+zzMO6y0t0zSmwGl0W4cNR5147hTSZjzMSYmyB61gmfHr2lA43i6VKhdKJg
XY6i+RBMwdQsjg+9084Abc8fr+fgPNAjZr8WhAPsHzPUVQdsaCK5hB3427fLnS6msAZRZ1sPx4CH
IOmSDcrzYpPGVRPTcyFLnJhovechBwHNZ1/nqm0NsR3k5W6M6RjMG/QIuZnu4rTLUt8uOu3udvQI
mAt9zBhwqE9PeXB9+qJnr34Bo4Kn+xk9ycjoilrFn+VJaYFqSwtLV2r011ACW4QB13IpWbMZk993
XIMw4bm/C8/OpPhULs6J3EONHRK0Wq9Q1r2TwiqgbXPIjhvS5yijM5ZOw9GvRoPz5TwXMuTHK+ty
MXvtocjf+vBbdxtNSe0wTmQeYKWYuHFmZtN+eZMEosHAZI+7mvod9FcXMHHHRfo+zbrYWKIKcIqe
X00cv0HCSHiBSV1vzNm6Adp//QKuKoWFunxUk6Z3PHbZ3DSzOE+akuNF7ZTVav0W0XGcw5Oj+m/F
aqITUMBcs7hdJfOxeMMDldU5/RLhI8NOkh2xTjF1sUfphPaPviWcBHAwp2hjSuNfYtHagiXyYx9x
muLIsUqLlhOgzWiJLNgesZyQ6QWPgT8hfC/pPtD1jYwDPWsX9WI8pqTau83fE3xLEJScBFU3Mv7I
0msKtb1GPMhApuNqRJ5l5Z+uNcL+0hH6Iw+/K2QhsZGiwT130lGZoQt+NfrOE+bryDCaPIKsNDXZ
WZPDkUJpol1a79iY5vq+Z7y6mOOQuvzmzujUfpOK0sjUdxtMzvqjrNn35AvDlPM9it1wI7aHoKZy
xbc/sVCWO1o+AcFlKgkZtVKDXMn1eL4xgVHtttuN/jrHqfdQ7t/RJk1dArdMpyNTNVFJuPcYnloR
6SUi6pUGAK25AA25m8e5fvPjCAHT+T9rvTnmXJ1emtE4MIFwVmiYVw9INmN48jASBfTB4Qncf8ov
XEq6If/W+JaMP5U7zkFfTiBFQysD04yMXdBxpWO/6iNOqnDlqDIsSqh2o8OrFDwJbyZ5rue3Ocjw
IyMmhQ6zb0Av1dnu8QvByhcCR/W+yme7OtghVoQ3GqXStanHQ9w14un90VqwdlGkn+ugEJKRWxJn
tLghKaUiCwa1wEP/w82KV24ITz1MFau/rmdsJznJUTUmF3xHGRmpmtIY/oqsaxyxY4e0LQYzz4kl
8W25GP1CD5ShxAZPmq8vLkB+yqZjfy0jkqkqRDpB69/4HeNi6p3vDNpqtljARwJ+IUC8Fk5fSMD9
7bWBod1VwgIzlFeh3zfRAunoh6PbzVQ1pxHuSZhDwJ+PRJD/uDZ1hDgI24SllkOLsnbsAA7M5Lsl
oCZFGsUD1RnAP2iB3BtZ6pp8EvBnP9Pqghs1ldKYyeJ9lwu+Q+q/fBeHcI86MgFV1rLsl8tcMo3+
uUX2OsyYTSWkG22Afe1RVkxMZvqSlbXRY2BkGH0hUmZHhSCiyd4q4MAkuOJQoVYDPFg5YHfvhkA5
/4Moy4LkYTfdMoWUpJstFu0ywgfegosqS5Wu4jphcVDoVB2b2McWUiE9LCjsTHkqpAfxejYNJFxu
GVs9vhhTNx8ya3LjadUrHbH3+SqffqDeKeHfbP8lc72P6bcVjEsaNQ/eI2jeXORhImf4SNM6lvob
iFwh/EWoUdVP7eQF6n4+FFqB4Ghi2llDF++Xy8r3iAv/EPjokeWH3ghvSJ6Z8ZPr4TMaF+xxau43
CYRlfWRr4tcq5NepV6UWBm8XKE+3JSjsIjY4fVFZblSg/EJDPAqQ/BS4mgOsyjxPAw5zoiAbkDeb
kXe4BAf+iHiAwmjyZjgJKZLNW03WpvhybsX5QUQp3kSo9Mq6wup9BuUzK23N6cpCZfAtSgZ37tIW
Pqn3xNrGodfItGAQTuHflOB+C56rcll20dqrrLtmPMSL+ieZn+B1ikfqhwOUVd965ji3CpQVu99P
ejoOzuq5uqY/qKciHLhcU8cv3UXRnBfEH66ll5UDOGOgkIa4qUseLEzj+d956WRUukIik1hZ48w5
U/rO5D63aDBIUt+hNg+N7SAgDwlmTlNACN0JPvAuIIs2AzsWXaYK772fgBuo59vQeMhOE/YSBNEq
X0vSsc3jht3/HybnW2YYyaIcW1JvzmIcF0ef7chyP8B2Du/fPG9syIOc0q4CBplF/7lUcM2TK3Ls
88LxI678ppOJO4fuappaDXIp3rSoOOpk7/kpKTQrtVxe+404R151+Gn5K96OQpl+cjC/T3QxVZHg
BE5msRTeU2f+zAJ2auaC0HDUndEsOsBlFSokIMskV9gJM9Wy5dyBG1sYJYmvwiYUGfoogWFl82mD
33o2nMlAjvt4TsFJ8lAPFD3ufHZ5mbWIfdhMF5rwNyJ3tHm214DbYo98KKmMi2nR5YqgmEb2fG38
jYhTjNq4YllbtfKfCPECYFw4nRbARYrPYuHqwisR3ByY6+MRSXwKtlcojALqvXROYAYI+0DFtvO0
GcV4Jl/uTjdXj2slk3EeAHW7hAxH9SBTjTDerEWoj6smxRbmZM+IKb7MSaVSaJX+EXUx87pClD+s
ge/w+8IH5RqF2Iac116SeeajXDxQYYla+4YoB+wJ6EgO1aThQJj/TDWR+rr5H1C7/BALJ9qHfXTW
Mj0DMAvZG2aeqFzzKrieBQOchf3PC8IvNiXCWZKqUyw1FeBiuynUmmxvxpshfSKYE1e2gmRoh2yi
KqaqipECtb4kL2+8OQ2EQZp6oOxJnhnjST8y4v/Vuqw0U7EkWUCpIszo/hoAos0ukLsafQcPzui4
5BwxbS9tivAtdTmDMeUSFXiAEUjQJQ9KjXe6M7BVdPvcSIpQWOWU/yF/6qb5Pq4MbhObdvm5A4IY
RYEdCe5naIVcI6w+tBBOHE7xwt5F7/mMsudzVCtJt6QGrOw/zXPYiWYbZSz3wCVrOOUNt5RnuQoE
p6f+6aSOdDUPy6FVqcqf9QlUQZsKm84ycSazO5sFtWzut7uzqeibamCnFz08xDIKnrCJsyG9ywSE
w8X8NKEPnNJ2P9vN0xVv/q4bAXVJpmalhIM/9FwdFo3sta7vTzWLj9L9siEJoY2Q3yy0JG4e2VDF
uiaj7WnxNkqKxZbGB1FwFFU9nrBTEdBgYLz//QdMiQ/c0Yk39uZVerCur8vK5gObdkIy32Vr77hK
lH0FZhOne4d6PsV7UpWF3saB62OQ/Bk8Y96KxsMZy6jot9XopAhpxLExWZUPy224DtVG5n+jvOOv
fLb+E8XlzIEa2d78sXhl7k897xlKr4NS/0G8p83NPytvuwv9XtU9bT5NTWHDj84hsFlZ3jYfgnHn
dwkOGw67ct1DKd2zEjlrY6Lmvf53H6KXskU6Mh0XlC8EqbIXOvDB/eHH2U8dYYOJJYp0is8t0gBw
6S000hdxVzHJ3VmUu9eidN5SH1+5PbeYUjVtr3T77f/2oi6jDZkuSzhnngsSxWSVJXzwZUQ6IYoW
7zW1HMpBn7sfhAdVX7IB7Nar+3iX0d9FaPadD8VGticdI02J77+lagAk2PIy2PIF3ErcTtvHkWDL
Lymz+QKfk20fgo1KRzE9iIDkN24xVxOcM3DuBTTSGWdCP9ikjFQqQjMO/ERzTwvHxwF0m7i73EFq
JW0VDCH7DjK+zlE6pVk2CVW71qneH3Z/nydkO8U3FZmlbPhCpHoQuqQ6vb/hjA9Wno4fIj+C+su7
F3AYepCtYJrcMuyHMab32hPfHSp6oZXO25btInVY2KeBTop07OR+de9BLp1peR8tDYTdeclJsZM9
KymIxGWDfKASUkVWnCinos/i/l71ZyRCT5UQSJx0KD3CQCZZj595l1A=
`protect end_protected

